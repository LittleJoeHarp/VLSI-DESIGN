magic
tech scmos
timestamp 1732047296
<< nwell >>
rect 4129 2122 4153 2146
rect 4339 2132 4390 2174
rect 4470 2143 4521 2169
rect 4553 2132 4604 2158
rect 4196 2107 4230 2113
rect 3326 2063 3377 2105
rect 3457 2074 3508 2100
rect 3540 2063 3591 2089
rect 3346 2021 3397 2055
rect 3620 2054 3658 2086
rect 4129 2067 4153 2091
rect 4168 2077 4230 2107
rect 4359 2090 4410 2124
rect 4633 2123 4671 2155
rect 4168 2071 4202 2077
rect 3765 1985 3789 2009
rect 3804 1999 3838 2005
rect 3804 1969 3866 1999
rect 3879 1970 3913 2006
rect 4021 2004 4055 2017
rect 4021 1981 4113 2004
rect 4055 1980 4113 1981
rect 3832 1963 3866 1969
rect 3333 1910 3384 1952
rect 3464 1921 3515 1947
rect 3547 1910 3598 1936
rect 3353 1868 3404 1902
rect 3627 1901 3665 1933
rect 3765 1930 3789 1954
rect 3929 1950 3963 1974
rect 4156 1948 4180 1972
rect 4223 1933 4257 1939
rect 4375 1933 4426 1975
rect 4506 1944 4557 1970
rect 4589 1933 4640 1959
rect 4156 1893 4180 1917
rect 4195 1903 4257 1933
rect 4195 1897 4229 1903
rect 4395 1891 4446 1925
rect 4669 1924 4707 1956
rect 3334 1759 3385 1801
rect 3465 1770 3516 1796
rect 3548 1759 3599 1785
rect 3354 1717 3405 1751
rect 3628 1750 3666 1782
rect 3765 1744 3789 1768
rect 3804 1758 3838 1764
rect 3804 1728 3866 1758
rect 3879 1729 3913 1765
rect 4016 1758 4050 1794
rect 4115 1761 4139 1762
rect 4081 1738 4139 1761
rect 4081 1737 4115 1738
rect 3832 1722 3866 1728
rect 3765 1689 3789 1713
rect 3929 1709 3963 1733
rect 4061 1707 4085 1731
rect 4095 1707 4129 1731
rect 4150 1725 4184 1738
rect 4150 1702 4208 1725
rect 4228 1702 4252 1726
rect 4267 1716 4301 1722
rect 4184 1701 4208 1702
rect 4016 1663 4050 1699
rect 4267 1686 4329 1716
rect 4295 1680 4329 1686
rect 4385 1680 4436 1722
rect 4516 1691 4567 1717
rect 4599 1680 4650 1706
rect 4228 1647 4252 1671
rect 3340 1604 3391 1646
rect 3471 1615 3522 1641
rect 4405 1638 4456 1672
rect 4679 1671 4717 1703
rect 3554 1604 3605 1630
rect 3360 1562 3411 1596
rect 3634 1595 3672 1627
rect 3765 1525 3789 1549
rect 3804 1539 3838 1545
rect 3804 1509 3866 1539
rect 3879 1510 3913 1546
rect 4016 1539 4050 1575
rect 4111 1542 4135 1543
rect 4077 1519 4135 1542
rect 4077 1518 4111 1519
rect 3832 1503 3866 1509
rect 3330 1457 3381 1499
rect 3461 1468 3512 1494
rect 3544 1457 3595 1483
rect 3350 1415 3401 1449
rect 3624 1448 3662 1480
rect 3765 1470 3789 1494
rect 3929 1490 3963 1514
rect 4061 1488 4085 1512
rect 4095 1488 4129 1512
rect 4149 1506 4183 1519
rect 4149 1483 4207 1506
rect 4225 1483 4249 1507
rect 4264 1497 4298 1503
rect 4183 1482 4207 1483
rect 4016 1444 4050 1480
rect 4264 1467 4326 1497
rect 4385 1467 4436 1509
rect 4516 1478 4567 1504
rect 4599 1467 4650 1493
rect 4292 1461 4326 1467
rect 4225 1428 4249 1452
rect 4405 1425 4456 1459
rect 4679 1458 4717 1490
rect 3331 1310 3382 1352
rect 3462 1321 3513 1347
rect 3545 1310 3596 1336
rect 3351 1268 3402 1302
rect 3625 1301 3663 1333
rect 3765 1302 3789 1326
rect 3804 1316 3838 1322
rect 3804 1286 3866 1316
rect 3879 1287 3913 1323
rect 4013 1316 4047 1352
rect 4254 1324 4278 1325
rect 4187 1323 4211 1324
rect 4109 1319 4133 1320
rect 4075 1296 4133 1319
rect 4153 1300 4211 1323
rect 4220 1301 4278 1324
rect 4220 1300 4254 1301
rect 4153 1299 4187 1300
rect 4075 1295 4109 1296
rect 3832 1280 3866 1286
rect 3765 1247 3789 1271
rect 3929 1267 3963 1291
rect 4058 1265 4082 1289
rect 4092 1265 4126 1289
rect 4140 1280 4174 1293
rect 4140 1257 4198 1280
rect 4013 1221 4047 1257
rect 4174 1256 4198 1257
rect 4207 1267 4241 1280
rect 4382 1277 4433 1319
rect 4513 1288 4564 1314
rect 4596 1277 4647 1303
rect 4207 1244 4265 1267
rect 4241 1243 4265 1244
rect 4402 1235 4453 1269
rect 4676 1268 4714 1300
rect 3340 1148 3391 1190
rect 3471 1159 3522 1185
rect 3554 1148 3605 1174
rect 3360 1106 3411 1140
rect 3634 1139 3672 1171
rect 3342 1010 3393 1052
rect 3473 1021 3524 1047
rect 3556 1010 3607 1036
rect 3362 968 3413 1002
rect 3636 1001 3674 1033
<< ntransistor >>
rect 4140 2154 4142 2160
rect 4179 2142 4181 2154
rect 4189 2142 4191 2154
rect 4207 2142 4209 2154
rect 4217 2142 4219 2154
rect 4140 2099 4142 2105
rect 4492 2107 4494 2119
rect 4579 2107 4581 2119
rect 4648 2087 4650 2093
rect 4381 2070 4383 2076
rect 4472 2075 4474 2087
rect 4555 2075 4557 2087
rect 3479 2038 3481 2050
rect 3566 2038 3568 2050
rect 3635 2018 3637 2024
rect 3368 2001 3370 2007
rect 3459 2006 3461 2018
rect 3542 2006 3544 2018
rect 3776 1971 3778 1977
rect 4066 1966 4068 1972
rect 4167 1980 4169 1986
rect 4206 1968 4208 1980
rect 4216 1968 4218 1980
rect 4234 1968 4236 1980
rect 4244 1968 4246 1980
rect 4032 1960 4034 1966
rect 4042 1960 4044 1966
rect 3890 1949 3892 1955
rect 3900 1949 3902 1955
rect 4090 1954 4092 1966
rect 4100 1954 4102 1966
rect 3815 1922 3817 1934
rect 3825 1922 3827 1934
rect 3843 1922 3845 1934
rect 3853 1922 3855 1934
rect 3940 1924 3942 1936
rect 3950 1924 3952 1936
rect 4167 1925 4169 1931
rect 3776 1916 3778 1922
rect 3486 1885 3488 1897
rect 3573 1885 3575 1897
rect 4528 1908 4530 1920
rect 4615 1908 4617 1920
rect 4684 1888 4686 1894
rect 4417 1871 4419 1877
rect 4508 1876 4510 1888
rect 4591 1876 4593 1888
rect 3642 1865 3644 1871
rect 3375 1848 3377 1854
rect 3466 1853 3468 1865
rect 3549 1853 3551 1865
rect 3487 1734 3489 1746
rect 3574 1734 3576 1746
rect 4092 1775 4094 1787
rect 4102 1775 4104 1787
rect 3776 1730 3778 1736
rect 4126 1770 4128 1776
rect 4027 1737 4029 1743
rect 4037 1737 4039 1743
rect 3643 1714 3645 1720
rect 3376 1697 3378 1703
rect 3467 1702 3469 1714
rect 3550 1702 3552 1714
rect 3890 1708 3892 1714
rect 3900 1708 3902 1714
rect 4027 1714 4029 1720
rect 4037 1714 4039 1720
rect 3815 1681 3817 1693
rect 3825 1681 3827 1693
rect 3843 1681 3845 1693
rect 3853 1681 3855 1693
rect 3940 1683 3942 1695
rect 3950 1683 3952 1695
rect 4072 1693 4074 1699
rect 3776 1675 3778 1681
rect 4106 1681 4108 1693
rect 4116 1681 4118 1693
rect 4195 1687 4197 1693
rect 4239 1688 4241 1694
rect 4161 1681 4163 1687
rect 4171 1681 4173 1687
rect 4278 1639 4280 1651
rect 4288 1639 4290 1651
rect 4306 1639 4308 1651
rect 4316 1639 4318 1651
rect 4239 1633 4241 1639
rect 4538 1655 4540 1667
rect 4625 1655 4627 1667
rect 4694 1635 4696 1641
rect 4427 1618 4429 1624
rect 4518 1623 4520 1635
rect 4601 1623 4603 1635
rect 3493 1579 3495 1591
rect 3580 1579 3582 1591
rect 3649 1559 3651 1565
rect 3382 1542 3384 1548
rect 3473 1547 3475 1559
rect 3556 1547 3558 1559
rect 4088 1556 4090 1568
rect 4098 1556 4100 1568
rect 3776 1511 3778 1517
rect 4122 1551 4124 1557
rect 4027 1518 4029 1524
rect 4037 1518 4039 1524
rect 3890 1489 3892 1495
rect 3900 1489 3902 1495
rect 4027 1495 4029 1501
rect 4037 1495 4039 1501
rect 3815 1462 3817 1474
rect 3825 1462 3827 1474
rect 3843 1462 3845 1474
rect 3853 1462 3855 1474
rect 3940 1464 3942 1476
rect 3950 1464 3952 1476
rect 4072 1474 4074 1480
rect 3483 1432 3485 1444
rect 3570 1432 3572 1444
rect 3776 1456 3778 1462
rect 4106 1462 4108 1474
rect 4116 1462 4118 1474
rect 4194 1468 4196 1474
rect 4236 1469 4238 1475
rect 4160 1462 4162 1468
rect 4170 1462 4172 1468
rect 4275 1420 4277 1432
rect 4285 1420 4287 1432
rect 4303 1420 4305 1432
rect 4313 1420 4315 1432
rect 3639 1412 3641 1418
rect 4236 1414 4238 1420
rect 4538 1442 4540 1454
rect 4625 1442 4627 1454
rect 4694 1422 4696 1428
rect 3372 1395 3374 1401
rect 3463 1400 3465 1412
rect 3546 1400 3548 1412
rect 4427 1405 4429 1411
rect 4518 1410 4520 1422
rect 4601 1410 4603 1422
rect 4086 1333 4088 1345
rect 4096 1333 4098 1345
rect 4164 1337 4166 1349
rect 4174 1337 4176 1349
rect 4231 1338 4233 1350
rect 4241 1338 4243 1350
rect 3484 1285 3486 1297
rect 3571 1285 3573 1297
rect 3776 1288 3778 1294
rect 4120 1328 4122 1334
rect 4198 1332 4200 1338
rect 4265 1333 4267 1339
rect 4024 1295 4026 1301
rect 4034 1295 4036 1301
rect 3640 1265 3642 1271
rect 3373 1248 3375 1254
rect 3464 1253 3466 1265
rect 3547 1253 3549 1265
rect 3890 1266 3892 1272
rect 3900 1266 3902 1272
rect 4024 1272 4026 1278
rect 4034 1272 4036 1278
rect 3815 1239 3817 1251
rect 3825 1239 3827 1251
rect 3843 1239 3845 1251
rect 3853 1239 3855 1251
rect 3940 1241 3942 1253
rect 3950 1241 3952 1253
rect 4069 1251 4071 1257
rect 3776 1233 3778 1239
rect 4103 1239 4105 1251
rect 4113 1239 4115 1251
rect 4185 1242 4187 1248
rect 4151 1236 4153 1242
rect 4161 1236 4163 1242
rect 4252 1229 4254 1235
rect 4218 1223 4220 1229
rect 4228 1223 4230 1229
rect 4535 1252 4537 1264
rect 4622 1252 4624 1264
rect 4691 1232 4693 1238
rect 4424 1215 4426 1221
rect 4515 1220 4517 1232
rect 4598 1220 4600 1232
rect 3493 1123 3495 1135
rect 3580 1123 3582 1135
rect 3649 1103 3651 1109
rect 3382 1086 3384 1092
rect 3473 1091 3475 1103
rect 3556 1091 3558 1103
rect 3495 985 3497 997
rect 3582 985 3584 997
rect 3651 965 3653 971
rect 3384 948 3386 954
rect 3475 953 3477 965
rect 3558 953 3560 965
<< ptransistor >>
rect 4140 2128 4142 2140
rect 4361 2139 4363 2163
rect 4492 2150 4494 2162
rect 3348 2070 3350 2094
rect 4575 2139 4577 2151
rect 3479 2081 3481 2093
rect 3562 2070 3564 2082
rect 3368 2027 3370 2049
rect 3635 2068 3637 2080
rect 4140 2073 4142 2085
rect 4179 2077 4181 2101
rect 4189 2077 4191 2101
rect 4207 2083 4209 2107
rect 4217 2083 4219 2107
rect 4381 2096 4383 2118
rect 4648 2137 4650 2149
rect 3776 1991 3778 2003
rect 3815 1975 3817 1999
rect 3825 1975 3827 1999
rect 3843 1969 3845 1993
rect 3853 1969 3855 1993
rect 3890 1976 3892 2000
rect 3900 1976 3902 2000
rect 4032 1987 4034 2011
rect 4042 1987 4044 2011
rect 3355 1917 3357 1941
rect 3486 1928 3488 1940
rect 3776 1936 3778 1948
rect 3569 1917 3571 1929
rect 3375 1874 3377 1896
rect 3642 1915 3644 1927
rect 3940 1956 3942 1968
rect 3950 1956 3952 1968
rect 4066 1986 4068 1998
rect 4090 1986 4092 1998
rect 4100 1986 4102 1998
rect 4167 1954 4169 1966
rect 4397 1940 4399 1964
rect 4528 1951 4530 1963
rect 4167 1899 4169 1911
rect 4206 1903 4208 1927
rect 4216 1903 4218 1927
rect 4234 1909 4236 1933
rect 4244 1909 4246 1933
rect 4611 1940 4613 1952
rect 4417 1897 4419 1919
rect 4684 1938 4686 1950
rect 3356 1766 3358 1790
rect 3487 1777 3489 1789
rect 3570 1766 3572 1778
rect 3376 1723 3378 1745
rect 3643 1764 3645 1776
rect 4027 1764 4029 1788
rect 4037 1764 4039 1788
rect 3776 1750 3778 1762
rect 3815 1734 3817 1758
rect 3825 1734 3827 1758
rect 3843 1728 3845 1752
rect 3853 1728 3855 1752
rect 3890 1735 3892 1759
rect 3900 1735 3902 1759
rect 4092 1743 4094 1755
rect 4102 1743 4104 1755
rect 4126 1744 4128 1756
rect 3776 1695 3778 1707
rect 3940 1715 3942 1727
rect 3950 1715 3952 1727
rect 4072 1713 4074 1725
rect 4106 1713 4108 1725
rect 4116 1713 4118 1725
rect 4161 1708 4163 1732
rect 4171 1708 4173 1732
rect 4027 1669 4029 1693
rect 4037 1669 4039 1693
rect 4195 1707 4197 1719
rect 4239 1708 4241 1720
rect 4278 1692 4280 1716
rect 4288 1692 4290 1716
rect 4306 1686 4308 1710
rect 4316 1686 4318 1710
rect 4407 1687 4409 1711
rect 4538 1698 4540 1710
rect 4239 1653 4241 1665
rect 3362 1611 3364 1635
rect 4621 1687 4623 1699
rect 3493 1622 3495 1634
rect 4427 1644 4429 1666
rect 4694 1685 4696 1697
rect 3576 1611 3578 1623
rect 3382 1568 3384 1590
rect 3649 1609 3651 1621
rect 4027 1545 4029 1569
rect 4037 1545 4039 1569
rect 3776 1531 3778 1543
rect 3815 1515 3817 1539
rect 3825 1515 3827 1539
rect 3843 1509 3845 1533
rect 3853 1509 3855 1533
rect 3890 1516 3892 1540
rect 3900 1516 3902 1540
rect 4088 1524 4090 1536
rect 4098 1524 4100 1536
rect 4122 1525 4124 1537
rect 3352 1464 3354 1488
rect 3483 1475 3485 1487
rect 3566 1464 3568 1476
rect 3776 1476 3778 1488
rect 3372 1421 3374 1443
rect 3639 1462 3641 1474
rect 3940 1496 3942 1508
rect 3950 1496 3952 1508
rect 4072 1494 4074 1506
rect 4106 1494 4108 1506
rect 4116 1494 4118 1506
rect 4160 1489 4162 1513
rect 4170 1489 4172 1513
rect 4027 1450 4029 1474
rect 4037 1450 4039 1474
rect 4194 1488 4196 1500
rect 4236 1489 4238 1501
rect 4275 1473 4277 1497
rect 4285 1473 4287 1497
rect 4303 1467 4305 1491
rect 4313 1467 4315 1491
rect 4407 1474 4409 1498
rect 4538 1485 4540 1497
rect 4236 1434 4238 1446
rect 4621 1474 4623 1486
rect 4427 1431 4429 1453
rect 4694 1472 4696 1484
rect 3353 1317 3355 1341
rect 3484 1328 3486 1340
rect 3567 1317 3569 1329
rect 3373 1274 3375 1296
rect 3640 1315 3642 1327
rect 4024 1322 4026 1346
rect 4034 1322 4036 1346
rect 3776 1308 3778 1320
rect 3815 1292 3817 1316
rect 3825 1292 3827 1316
rect 3843 1286 3845 1310
rect 3853 1286 3855 1310
rect 3890 1293 3892 1317
rect 3900 1293 3902 1317
rect 4086 1301 4088 1313
rect 4096 1301 4098 1313
rect 4120 1302 4122 1314
rect 4164 1305 4166 1317
rect 4174 1305 4176 1317
rect 4198 1306 4200 1318
rect 4231 1306 4233 1318
rect 4241 1306 4243 1318
rect 4265 1307 4267 1319
rect 3776 1253 3778 1265
rect 3940 1273 3942 1285
rect 3950 1273 3952 1285
rect 4069 1271 4071 1283
rect 4103 1271 4105 1283
rect 4113 1271 4115 1283
rect 4151 1263 4153 1287
rect 4161 1263 4163 1287
rect 4404 1284 4406 1308
rect 4535 1295 4537 1307
rect 4024 1227 4026 1251
rect 4034 1227 4036 1251
rect 4185 1262 4187 1274
rect 4218 1250 4220 1274
rect 4228 1250 4230 1274
rect 4618 1284 4620 1296
rect 4252 1249 4254 1261
rect 4424 1241 4426 1263
rect 4691 1282 4693 1294
rect 3362 1155 3364 1179
rect 3493 1166 3495 1178
rect 3576 1155 3578 1167
rect 3382 1112 3384 1134
rect 3649 1153 3651 1165
rect 3364 1017 3366 1041
rect 3495 1028 3497 1040
rect 3578 1017 3580 1029
rect 3384 974 3386 996
rect 3651 1015 3653 1027
<< ndiffusion >>
rect 4139 2154 4140 2160
rect 4142 2154 4143 2160
rect 4178 2142 4179 2154
rect 4181 2142 4189 2154
rect 4191 2142 4192 2154
rect 4206 2142 4207 2154
rect 4209 2142 4217 2154
rect 4219 2142 4220 2154
rect 4139 2099 4140 2105
rect 4142 2099 4143 2105
rect 4478 2112 4492 2119
rect 4478 2107 4480 2112
rect 4489 2107 4492 2112
rect 4494 2113 4500 2119
rect 4509 2113 4519 2119
rect 4494 2107 4519 2113
rect 4559 2112 4579 2119
rect 4559 2107 4561 2112
rect 4570 2107 4579 2112
rect 4581 2113 4583 2119
rect 4592 2113 4602 2119
rect 4581 2107 4602 2113
rect 4638 2091 4648 2093
rect 4638 2087 4639 2091
rect 4646 2087 4648 2091
rect 4650 2087 4653 2093
rect 4664 2087 4677 2093
rect 4458 2080 4472 2087
rect 4367 2075 4381 2076
rect 4367 2070 4369 2075
rect 4377 2070 4381 2075
rect 4383 2070 4389 2076
rect 4398 2070 4408 2076
rect 4458 2075 4460 2080
rect 4468 2075 4472 2080
rect 4474 2081 4480 2087
rect 4489 2081 4499 2087
rect 4474 2075 4499 2081
rect 4541 2080 4555 2087
rect 4541 2075 4543 2080
rect 4551 2075 4555 2080
rect 4557 2081 4561 2087
rect 4570 2081 4582 2087
rect 4557 2075 4582 2081
rect 3465 2043 3479 2050
rect 3465 2038 3467 2043
rect 3476 2038 3479 2043
rect 3481 2044 3487 2050
rect 3496 2044 3506 2050
rect 3481 2038 3506 2044
rect 3546 2043 3566 2050
rect 3546 2038 3548 2043
rect 3557 2038 3566 2043
rect 3568 2044 3570 2050
rect 3579 2044 3589 2050
rect 3568 2038 3589 2044
rect 3625 2022 3635 2024
rect 3625 2018 3626 2022
rect 3633 2018 3635 2022
rect 3637 2018 3640 2024
rect 3651 2018 3664 2024
rect 3445 2011 3459 2018
rect 3354 2006 3368 2007
rect 3354 2001 3356 2006
rect 3364 2001 3368 2006
rect 3370 2001 3376 2007
rect 3385 2001 3395 2007
rect 3445 2006 3447 2011
rect 3455 2006 3459 2011
rect 3461 2012 3467 2018
rect 3476 2012 3486 2018
rect 3461 2006 3486 2012
rect 3528 2011 3542 2018
rect 3528 2006 3530 2011
rect 3538 2006 3542 2011
rect 3544 2012 3548 2018
rect 3557 2012 3569 2018
rect 3544 2006 3569 2012
rect 3775 1971 3776 1977
rect 3778 1971 3779 1977
rect 4065 1966 4066 1972
rect 4068 1966 4069 1972
rect 4166 1980 4167 1986
rect 4169 1980 4170 1986
rect 4205 1968 4206 1980
rect 4208 1968 4216 1980
rect 4218 1968 4219 1980
rect 4233 1968 4234 1980
rect 4236 1968 4244 1980
rect 4246 1968 4247 1980
rect 4031 1960 4032 1966
rect 4034 1960 4036 1966
rect 4040 1960 4042 1966
rect 4044 1960 4045 1966
rect 3889 1949 3890 1955
rect 3892 1949 3894 1955
rect 3898 1949 3900 1955
rect 3902 1949 3903 1955
rect 4089 1954 4090 1966
rect 4092 1954 4100 1966
rect 4102 1954 4103 1966
rect 3814 1922 3815 1934
rect 3817 1922 3825 1934
rect 3827 1922 3828 1934
rect 3842 1922 3843 1934
rect 3845 1922 3853 1934
rect 3855 1922 3856 1934
rect 3939 1924 3940 1936
rect 3942 1924 3950 1936
rect 3952 1924 3953 1936
rect 4166 1925 4167 1931
rect 4169 1925 4170 1931
rect 3775 1916 3776 1922
rect 3778 1916 3779 1922
rect 3472 1890 3486 1897
rect 3472 1885 3474 1890
rect 3483 1885 3486 1890
rect 3488 1891 3494 1897
rect 3503 1891 3513 1897
rect 3488 1885 3513 1891
rect 3553 1890 3573 1897
rect 3553 1885 3555 1890
rect 3564 1885 3573 1890
rect 3575 1891 3577 1897
rect 3586 1891 3596 1897
rect 3575 1885 3596 1891
rect 4514 1913 4528 1920
rect 4514 1908 4516 1913
rect 4525 1908 4528 1913
rect 4530 1914 4536 1920
rect 4545 1914 4555 1920
rect 4530 1908 4555 1914
rect 4595 1913 4615 1920
rect 4595 1908 4597 1913
rect 4606 1908 4615 1913
rect 4617 1914 4619 1920
rect 4628 1914 4638 1920
rect 4617 1908 4638 1914
rect 4674 1892 4684 1894
rect 4674 1888 4675 1892
rect 4682 1888 4684 1892
rect 4686 1888 4689 1894
rect 4700 1888 4713 1894
rect 4494 1881 4508 1888
rect 4403 1876 4417 1877
rect 4403 1871 4405 1876
rect 4413 1871 4417 1876
rect 4419 1871 4425 1877
rect 4434 1871 4444 1877
rect 4494 1876 4496 1881
rect 4504 1876 4508 1881
rect 4510 1882 4516 1888
rect 4525 1882 4535 1888
rect 4510 1876 4535 1882
rect 4577 1881 4591 1888
rect 4577 1876 4579 1881
rect 4587 1876 4591 1881
rect 4593 1882 4597 1888
rect 4606 1882 4618 1888
rect 4593 1876 4618 1882
rect 3632 1869 3642 1871
rect 3632 1865 3633 1869
rect 3640 1865 3642 1869
rect 3644 1865 3647 1871
rect 3658 1865 3671 1871
rect 3452 1858 3466 1865
rect 3361 1853 3375 1854
rect 3361 1848 3363 1853
rect 3371 1848 3375 1853
rect 3377 1848 3383 1854
rect 3392 1848 3402 1854
rect 3452 1853 3454 1858
rect 3462 1853 3466 1858
rect 3468 1859 3474 1865
rect 3483 1859 3493 1865
rect 3468 1853 3493 1859
rect 3535 1858 3549 1865
rect 3535 1853 3537 1858
rect 3545 1853 3549 1858
rect 3551 1859 3555 1865
rect 3564 1859 3576 1865
rect 3551 1853 3576 1859
rect 3473 1739 3487 1746
rect 3473 1734 3475 1739
rect 3484 1734 3487 1739
rect 3489 1740 3495 1746
rect 3504 1740 3514 1746
rect 3489 1734 3514 1740
rect 3554 1739 3574 1746
rect 3554 1734 3556 1739
rect 3565 1734 3574 1739
rect 3576 1740 3578 1746
rect 3587 1740 3597 1746
rect 3576 1734 3597 1740
rect 4091 1775 4092 1787
rect 4094 1775 4102 1787
rect 4104 1775 4105 1787
rect 3775 1730 3776 1736
rect 3778 1730 3779 1736
rect 4125 1770 4126 1776
rect 4128 1770 4129 1776
rect 4026 1737 4027 1743
rect 4029 1737 4031 1743
rect 4035 1737 4037 1743
rect 4039 1737 4040 1743
rect 3633 1718 3643 1720
rect 3633 1714 3634 1718
rect 3641 1714 3643 1718
rect 3645 1714 3648 1720
rect 3659 1714 3672 1720
rect 3453 1707 3467 1714
rect 3362 1702 3376 1703
rect 3362 1697 3364 1702
rect 3372 1697 3376 1702
rect 3378 1697 3384 1703
rect 3393 1697 3403 1703
rect 3453 1702 3455 1707
rect 3463 1702 3467 1707
rect 3469 1708 3475 1714
rect 3484 1708 3494 1714
rect 3469 1702 3494 1708
rect 3536 1707 3550 1714
rect 3536 1702 3538 1707
rect 3546 1702 3550 1707
rect 3552 1708 3556 1714
rect 3565 1708 3577 1714
rect 3552 1702 3577 1708
rect 3889 1708 3890 1714
rect 3892 1708 3894 1714
rect 3898 1708 3900 1714
rect 3902 1708 3903 1714
rect 4026 1714 4027 1720
rect 4029 1714 4031 1720
rect 4035 1714 4037 1720
rect 4039 1714 4040 1720
rect 3814 1681 3815 1693
rect 3817 1681 3825 1693
rect 3827 1681 3828 1693
rect 3842 1681 3843 1693
rect 3845 1681 3853 1693
rect 3855 1681 3856 1693
rect 3939 1683 3940 1695
rect 3942 1683 3950 1695
rect 3952 1683 3953 1695
rect 4071 1693 4072 1699
rect 4074 1693 4075 1699
rect 3775 1675 3776 1681
rect 3778 1675 3779 1681
rect 4105 1681 4106 1693
rect 4108 1681 4116 1693
rect 4118 1681 4119 1693
rect 4194 1687 4195 1693
rect 4197 1687 4198 1693
rect 4238 1688 4239 1694
rect 4241 1688 4242 1694
rect 4160 1681 4161 1687
rect 4163 1681 4165 1687
rect 4169 1681 4171 1687
rect 4173 1681 4174 1687
rect 4277 1639 4278 1651
rect 4280 1639 4288 1651
rect 4290 1639 4291 1651
rect 4305 1639 4306 1651
rect 4308 1639 4316 1651
rect 4318 1639 4319 1651
rect 4238 1633 4239 1639
rect 4241 1633 4242 1639
rect 4524 1660 4538 1667
rect 4524 1655 4526 1660
rect 4535 1655 4538 1660
rect 4540 1661 4546 1667
rect 4555 1661 4565 1667
rect 4540 1655 4565 1661
rect 4605 1660 4625 1667
rect 4605 1655 4607 1660
rect 4616 1655 4625 1660
rect 4627 1661 4629 1667
rect 4638 1661 4648 1667
rect 4627 1655 4648 1661
rect 4684 1639 4694 1641
rect 4684 1635 4685 1639
rect 4692 1635 4694 1639
rect 4696 1635 4699 1641
rect 4710 1635 4723 1641
rect 4504 1628 4518 1635
rect 4413 1623 4427 1624
rect 4413 1618 4415 1623
rect 4423 1618 4427 1623
rect 4429 1618 4435 1624
rect 4444 1618 4454 1624
rect 4504 1623 4506 1628
rect 4514 1623 4518 1628
rect 4520 1629 4526 1635
rect 4535 1629 4545 1635
rect 4520 1623 4545 1629
rect 4587 1628 4601 1635
rect 4587 1623 4589 1628
rect 4597 1623 4601 1628
rect 4603 1629 4607 1635
rect 4616 1629 4628 1635
rect 4603 1623 4628 1629
rect 3479 1584 3493 1591
rect 3479 1579 3481 1584
rect 3490 1579 3493 1584
rect 3495 1585 3501 1591
rect 3510 1585 3520 1591
rect 3495 1579 3520 1585
rect 3560 1584 3580 1591
rect 3560 1579 3562 1584
rect 3571 1579 3580 1584
rect 3582 1585 3584 1591
rect 3593 1585 3603 1591
rect 3582 1579 3603 1585
rect 3639 1563 3649 1565
rect 3639 1559 3640 1563
rect 3647 1559 3649 1563
rect 3651 1559 3654 1565
rect 3665 1559 3678 1565
rect 3459 1552 3473 1559
rect 3368 1547 3382 1548
rect 3368 1542 3370 1547
rect 3378 1542 3382 1547
rect 3384 1542 3390 1548
rect 3399 1542 3409 1548
rect 3459 1547 3461 1552
rect 3469 1547 3473 1552
rect 3475 1553 3481 1559
rect 3490 1553 3500 1559
rect 3475 1547 3500 1553
rect 3542 1552 3556 1559
rect 3542 1547 3544 1552
rect 3552 1547 3556 1552
rect 3558 1553 3562 1559
rect 3571 1553 3583 1559
rect 3558 1547 3583 1553
rect 4087 1556 4088 1568
rect 4090 1556 4098 1568
rect 4100 1556 4101 1568
rect 3775 1511 3776 1517
rect 3778 1511 3779 1517
rect 4121 1551 4122 1557
rect 4124 1551 4125 1557
rect 4026 1518 4027 1524
rect 4029 1518 4031 1524
rect 4035 1518 4037 1524
rect 4039 1518 4040 1524
rect 3889 1489 3890 1495
rect 3892 1489 3894 1495
rect 3898 1489 3900 1495
rect 3902 1489 3903 1495
rect 4026 1495 4027 1501
rect 4029 1495 4031 1501
rect 4035 1495 4037 1501
rect 4039 1495 4040 1501
rect 3814 1462 3815 1474
rect 3817 1462 3825 1474
rect 3827 1462 3828 1474
rect 3842 1462 3843 1474
rect 3845 1462 3853 1474
rect 3855 1462 3856 1474
rect 3939 1464 3940 1476
rect 3942 1464 3950 1476
rect 3952 1464 3953 1476
rect 4071 1474 4072 1480
rect 4074 1474 4075 1480
rect 3469 1437 3483 1444
rect 3469 1432 3471 1437
rect 3480 1432 3483 1437
rect 3485 1438 3491 1444
rect 3500 1438 3510 1444
rect 3485 1432 3510 1438
rect 3550 1437 3570 1444
rect 3550 1432 3552 1437
rect 3561 1432 3570 1437
rect 3572 1438 3574 1444
rect 3583 1438 3593 1444
rect 3572 1432 3593 1438
rect 3775 1456 3776 1462
rect 3778 1456 3779 1462
rect 4105 1462 4106 1474
rect 4108 1462 4116 1474
rect 4118 1462 4119 1474
rect 4193 1468 4194 1474
rect 4196 1468 4197 1474
rect 4235 1469 4236 1475
rect 4238 1469 4239 1475
rect 4159 1462 4160 1468
rect 4162 1462 4164 1468
rect 4168 1462 4170 1468
rect 4172 1462 4173 1468
rect 4274 1420 4275 1432
rect 4277 1420 4285 1432
rect 4287 1420 4288 1432
rect 4302 1420 4303 1432
rect 4305 1420 4313 1432
rect 4315 1420 4316 1432
rect 3629 1416 3639 1418
rect 3629 1412 3630 1416
rect 3637 1412 3639 1416
rect 3641 1412 3644 1418
rect 3655 1412 3668 1418
rect 4235 1414 4236 1420
rect 4238 1414 4239 1420
rect 4524 1447 4538 1454
rect 4524 1442 4526 1447
rect 4535 1442 4538 1447
rect 4540 1448 4546 1454
rect 4555 1448 4565 1454
rect 4540 1442 4565 1448
rect 4605 1447 4625 1454
rect 4605 1442 4607 1447
rect 4616 1442 4625 1447
rect 4627 1448 4629 1454
rect 4638 1448 4648 1454
rect 4627 1442 4648 1448
rect 4684 1426 4694 1428
rect 4684 1422 4685 1426
rect 4692 1422 4694 1426
rect 4696 1422 4699 1428
rect 4710 1422 4723 1428
rect 4504 1415 4518 1422
rect 3449 1405 3463 1412
rect 3358 1400 3372 1401
rect 3358 1395 3360 1400
rect 3368 1395 3372 1400
rect 3374 1395 3380 1401
rect 3389 1395 3399 1401
rect 3449 1400 3451 1405
rect 3459 1400 3463 1405
rect 3465 1406 3471 1412
rect 3480 1406 3490 1412
rect 3465 1400 3490 1406
rect 3532 1405 3546 1412
rect 3532 1400 3534 1405
rect 3542 1400 3546 1405
rect 3548 1406 3552 1412
rect 3561 1406 3573 1412
rect 3548 1400 3573 1406
rect 4413 1410 4427 1411
rect 4413 1405 4415 1410
rect 4423 1405 4427 1410
rect 4429 1405 4435 1411
rect 4444 1405 4454 1411
rect 4504 1410 4506 1415
rect 4514 1410 4518 1415
rect 4520 1416 4526 1422
rect 4535 1416 4545 1422
rect 4520 1410 4545 1416
rect 4587 1415 4601 1422
rect 4587 1410 4589 1415
rect 4597 1410 4601 1415
rect 4603 1416 4607 1422
rect 4616 1416 4628 1422
rect 4603 1410 4628 1416
rect 4085 1333 4086 1345
rect 4088 1333 4096 1345
rect 4098 1333 4099 1345
rect 4163 1337 4164 1349
rect 4166 1337 4174 1349
rect 4176 1337 4177 1349
rect 4230 1338 4231 1350
rect 4233 1338 4241 1350
rect 4243 1338 4244 1350
rect 3470 1290 3484 1297
rect 3470 1285 3472 1290
rect 3481 1285 3484 1290
rect 3486 1291 3492 1297
rect 3501 1291 3511 1297
rect 3486 1285 3511 1291
rect 3551 1290 3571 1297
rect 3551 1285 3553 1290
rect 3562 1285 3571 1290
rect 3573 1291 3575 1297
rect 3584 1291 3594 1297
rect 3573 1285 3594 1291
rect 3775 1288 3776 1294
rect 3778 1288 3779 1294
rect 4119 1328 4120 1334
rect 4122 1328 4123 1334
rect 4197 1332 4198 1338
rect 4200 1332 4201 1338
rect 4264 1333 4265 1339
rect 4267 1333 4268 1339
rect 4023 1295 4024 1301
rect 4026 1295 4028 1301
rect 4032 1295 4034 1301
rect 4036 1295 4037 1301
rect 3630 1269 3640 1271
rect 3630 1265 3631 1269
rect 3638 1265 3640 1269
rect 3642 1265 3645 1271
rect 3656 1265 3669 1271
rect 3450 1258 3464 1265
rect 3359 1253 3373 1254
rect 3359 1248 3361 1253
rect 3369 1248 3373 1253
rect 3375 1248 3381 1254
rect 3390 1248 3400 1254
rect 3450 1253 3452 1258
rect 3460 1253 3464 1258
rect 3466 1259 3472 1265
rect 3481 1259 3491 1265
rect 3466 1253 3491 1259
rect 3533 1258 3547 1265
rect 3533 1253 3535 1258
rect 3543 1253 3547 1258
rect 3549 1259 3553 1265
rect 3562 1259 3574 1265
rect 3549 1253 3574 1259
rect 3889 1266 3890 1272
rect 3892 1266 3894 1272
rect 3898 1266 3900 1272
rect 3902 1266 3903 1272
rect 4023 1272 4024 1278
rect 4026 1272 4028 1278
rect 4032 1272 4034 1278
rect 4036 1272 4037 1278
rect 3814 1239 3815 1251
rect 3817 1239 3825 1251
rect 3827 1239 3828 1251
rect 3842 1239 3843 1251
rect 3845 1239 3853 1251
rect 3855 1239 3856 1251
rect 3939 1241 3940 1253
rect 3942 1241 3950 1253
rect 3952 1241 3953 1253
rect 4068 1251 4069 1257
rect 4071 1251 4072 1257
rect 3775 1233 3776 1239
rect 3778 1233 3779 1239
rect 4102 1239 4103 1251
rect 4105 1239 4113 1251
rect 4115 1239 4116 1251
rect 4184 1242 4185 1248
rect 4187 1242 4188 1248
rect 4150 1236 4151 1242
rect 4153 1236 4155 1242
rect 4159 1236 4161 1242
rect 4163 1236 4164 1242
rect 4251 1229 4252 1235
rect 4254 1229 4255 1235
rect 4217 1223 4218 1229
rect 4220 1223 4222 1229
rect 4226 1223 4228 1229
rect 4230 1223 4231 1229
rect 4521 1257 4535 1264
rect 4521 1252 4523 1257
rect 4532 1252 4535 1257
rect 4537 1258 4543 1264
rect 4552 1258 4562 1264
rect 4537 1252 4562 1258
rect 4602 1257 4622 1264
rect 4602 1252 4604 1257
rect 4613 1252 4622 1257
rect 4624 1258 4626 1264
rect 4635 1258 4645 1264
rect 4624 1252 4645 1258
rect 4681 1236 4691 1238
rect 4681 1232 4682 1236
rect 4689 1232 4691 1236
rect 4693 1232 4696 1238
rect 4707 1232 4720 1238
rect 4501 1225 4515 1232
rect 4410 1220 4424 1221
rect 4410 1215 4412 1220
rect 4420 1215 4424 1220
rect 4426 1215 4432 1221
rect 4441 1215 4451 1221
rect 4501 1220 4503 1225
rect 4511 1220 4515 1225
rect 4517 1226 4523 1232
rect 4532 1226 4542 1232
rect 4517 1220 4542 1226
rect 4584 1225 4598 1232
rect 4584 1220 4586 1225
rect 4594 1220 4598 1225
rect 4600 1226 4604 1232
rect 4613 1226 4625 1232
rect 4600 1220 4625 1226
rect 3479 1128 3493 1135
rect 3479 1123 3481 1128
rect 3490 1123 3493 1128
rect 3495 1129 3501 1135
rect 3510 1129 3520 1135
rect 3495 1123 3520 1129
rect 3560 1128 3580 1135
rect 3560 1123 3562 1128
rect 3571 1123 3580 1128
rect 3582 1129 3584 1135
rect 3593 1129 3603 1135
rect 3582 1123 3603 1129
rect 3639 1107 3649 1109
rect 3639 1103 3640 1107
rect 3647 1103 3649 1107
rect 3651 1103 3654 1109
rect 3665 1103 3678 1109
rect 3459 1096 3473 1103
rect 3368 1091 3382 1092
rect 3368 1086 3370 1091
rect 3378 1086 3382 1091
rect 3384 1086 3390 1092
rect 3399 1086 3409 1092
rect 3459 1091 3461 1096
rect 3469 1091 3473 1096
rect 3475 1097 3481 1103
rect 3490 1097 3500 1103
rect 3475 1091 3500 1097
rect 3542 1096 3556 1103
rect 3542 1091 3544 1096
rect 3552 1091 3556 1096
rect 3558 1097 3562 1103
rect 3571 1097 3583 1103
rect 3558 1091 3583 1097
rect 3481 990 3495 997
rect 3481 985 3483 990
rect 3492 985 3495 990
rect 3497 991 3503 997
rect 3512 991 3522 997
rect 3497 985 3522 991
rect 3562 990 3582 997
rect 3562 985 3564 990
rect 3573 985 3582 990
rect 3584 991 3586 997
rect 3595 991 3605 997
rect 3584 985 3605 991
rect 3641 969 3651 971
rect 3641 965 3642 969
rect 3649 965 3651 969
rect 3653 965 3656 971
rect 3667 965 3680 971
rect 3461 958 3475 965
rect 3370 953 3384 954
rect 3370 948 3372 953
rect 3380 948 3384 953
rect 3386 948 3392 954
rect 3401 948 3411 954
rect 3461 953 3463 958
rect 3471 953 3475 958
rect 3477 959 3483 965
rect 3492 959 3502 965
rect 3477 953 3502 959
rect 3544 958 3558 965
rect 3544 953 3546 958
rect 3554 953 3558 958
rect 3560 959 3564 965
rect 3573 959 3585 965
rect 3560 953 3585 959
<< pdiffusion >>
rect 4346 2151 4361 2163
rect 4346 2142 4349 2151
rect 4357 2142 4361 2151
rect 4139 2128 4140 2140
rect 4142 2128 4143 2140
rect 4346 2139 4361 2142
rect 4363 2143 4381 2163
rect 4477 2153 4480 2162
rect 4488 2153 4492 2162
rect 4477 2150 4492 2153
rect 4494 2154 4512 2162
rect 4494 2150 4500 2154
rect 4509 2150 4512 2154
rect 4363 2139 4369 2143
rect 4378 2139 4381 2143
rect 4560 2142 4563 2151
rect 4571 2142 4575 2151
rect 3333 2082 3348 2094
rect 3333 2073 3336 2082
rect 3344 2073 3348 2082
rect 3333 2070 3348 2073
rect 3350 2074 3368 2094
rect 4560 2139 4575 2142
rect 4577 2143 4595 2151
rect 4577 2139 4583 2143
rect 4592 2139 4595 2143
rect 4639 2142 4640 2149
rect 4646 2142 4648 2149
rect 3464 2084 3467 2093
rect 3475 2084 3479 2093
rect 3464 2081 3479 2084
rect 3481 2085 3499 2093
rect 3481 2081 3487 2085
rect 3496 2081 3499 2085
rect 3350 2070 3356 2074
rect 3365 2070 3368 2074
rect 3547 2073 3550 2082
rect 3558 2073 3562 2082
rect 3547 2070 3562 2073
rect 3564 2074 3582 2082
rect 3564 2070 3570 2074
rect 3579 2070 3582 2074
rect 3626 2073 3627 2080
rect 3633 2073 3635 2080
rect 3353 2043 3368 2049
rect 3353 2034 3356 2043
rect 3365 2034 3368 2043
rect 3353 2027 3368 2034
rect 3370 2035 3388 2049
rect 3370 2031 3376 2035
rect 3385 2031 3388 2035
rect 3370 2027 3388 2031
rect 3626 2068 3635 2073
rect 3637 2073 3652 2080
rect 4139 2073 4140 2085
rect 4142 2073 4143 2085
rect 4178 2077 4179 2101
rect 4181 2077 4183 2101
rect 4187 2077 4189 2101
rect 4191 2077 4192 2101
rect 4206 2083 4207 2107
rect 4209 2083 4211 2107
rect 4215 2083 4217 2107
rect 4219 2083 4220 2107
rect 4366 2112 4381 2118
rect 4366 2103 4369 2112
rect 4378 2103 4381 2112
rect 4366 2096 4381 2103
rect 4383 2104 4401 2118
rect 4383 2100 4389 2104
rect 4398 2100 4401 2104
rect 4383 2096 4401 2100
rect 4639 2137 4648 2142
rect 4650 2142 4665 2149
rect 4650 2137 4653 2142
rect 4664 2137 4665 2142
rect 3637 2068 3640 2073
rect 3651 2068 3652 2073
rect 3775 1991 3776 2003
rect 3778 1991 3779 2003
rect 3814 1975 3815 1999
rect 3817 1975 3819 1999
rect 3823 1975 3825 1999
rect 3827 1975 3828 1999
rect 3842 1969 3843 1993
rect 3845 1969 3847 1993
rect 3851 1969 3853 1993
rect 3855 1969 3856 1993
rect 3889 1976 3890 2000
rect 3892 1976 3900 2000
rect 3902 1976 3903 2000
rect 4031 1987 4032 2011
rect 4034 1987 4042 2011
rect 4044 1987 4045 2011
rect 3340 1929 3355 1941
rect 3340 1920 3343 1929
rect 3351 1920 3355 1929
rect 3340 1917 3355 1920
rect 3357 1921 3375 1941
rect 3471 1931 3474 1940
rect 3482 1931 3486 1940
rect 3471 1928 3486 1931
rect 3488 1932 3506 1940
rect 3775 1936 3776 1948
rect 3778 1936 3779 1948
rect 3488 1928 3494 1932
rect 3503 1928 3506 1932
rect 3357 1917 3363 1921
rect 3372 1917 3375 1921
rect 3554 1920 3557 1929
rect 3565 1920 3569 1929
rect 3554 1917 3569 1920
rect 3571 1921 3589 1929
rect 3571 1917 3577 1921
rect 3586 1917 3589 1921
rect 3633 1920 3634 1927
rect 3640 1920 3642 1927
rect 3360 1890 3375 1896
rect 3360 1881 3363 1890
rect 3372 1881 3375 1890
rect 3360 1874 3375 1881
rect 3377 1882 3395 1896
rect 3377 1878 3383 1882
rect 3392 1878 3395 1882
rect 3377 1874 3395 1878
rect 3633 1915 3642 1920
rect 3644 1920 3659 1927
rect 3939 1956 3940 1968
rect 3942 1956 3944 1968
rect 3948 1956 3950 1968
rect 3952 1956 3953 1968
rect 4065 1986 4066 1998
rect 4068 1986 4069 1998
rect 4089 1986 4090 1998
rect 4092 1986 4094 1998
rect 4098 1986 4100 1998
rect 4102 1986 4103 1998
rect 4166 1954 4167 1966
rect 4169 1954 4170 1966
rect 4382 1952 4397 1964
rect 4382 1943 4385 1952
rect 4393 1943 4397 1952
rect 4382 1940 4397 1943
rect 4399 1944 4417 1964
rect 4513 1954 4516 1963
rect 4524 1954 4528 1963
rect 4513 1951 4528 1954
rect 4530 1955 4548 1963
rect 4530 1951 4536 1955
rect 4545 1951 4548 1955
rect 4399 1940 4405 1944
rect 4414 1940 4417 1944
rect 4596 1943 4599 1952
rect 4607 1943 4611 1952
rect 3644 1915 3647 1920
rect 3658 1915 3659 1920
rect 4166 1899 4167 1911
rect 4169 1899 4170 1911
rect 4205 1903 4206 1927
rect 4208 1903 4210 1927
rect 4214 1903 4216 1927
rect 4218 1903 4219 1927
rect 4233 1909 4234 1933
rect 4236 1909 4238 1933
rect 4242 1909 4244 1933
rect 4246 1909 4247 1933
rect 4596 1940 4611 1943
rect 4613 1944 4631 1952
rect 4613 1940 4619 1944
rect 4628 1940 4631 1944
rect 4675 1943 4676 1950
rect 4682 1943 4684 1950
rect 4402 1913 4417 1919
rect 4402 1904 4405 1913
rect 4414 1904 4417 1913
rect 4402 1897 4417 1904
rect 4419 1905 4437 1919
rect 4419 1901 4425 1905
rect 4434 1901 4437 1905
rect 4419 1897 4437 1901
rect 4675 1938 4684 1943
rect 4686 1943 4701 1950
rect 4686 1938 4689 1943
rect 4700 1938 4701 1943
rect 3341 1778 3356 1790
rect 3341 1769 3344 1778
rect 3352 1769 3356 1778
rect 3341 1766 3356 1769
rect 3358 1770 3376 1790
rect 3472 1780 3475 1789
rect 3483 1780 3487 1789
rect 3472 1777 3487 1780
rect 3489 1781 3507 1789
rect 3489 1777 3495 1781
rect 3504 1777 3507 1781
rect 3358 1766 3364 1770
rect 3373 1766 3376 1770
rect 3555 1769 3558 1778
rect 3566 1769 3570 1778
rect 3555 1766 3570 1769
rect 3572 1770 3590 1778
rect 3572 1766 3578 1770
rect 3587 1766 3590 1770
rect 3634 1769 3635 1776
rect 3641 1769 3643 1776
rect 3361 1739 3376 1745
rect 3361 1730 3364 1739
rect 3373 1730 3376 1739
rect 3361 1723 3376 1730
rect 3378 1731 3396 1745
rect 3378 1727 3384 1731
rect 3393 1727 3396 1731
rect 3378 1723 3396 1727
rect 3634 1764 3643 1769
rect 3645 1769 3660 1776
rect 3645 1764 3648 1769
rect 3659 1764 3660 1769
rect 4026 1764 4027 1788
rect 4029 1764 4037 1788
rect 4039 1764 4040 1788
rect 3775 1750 3776 1762
rect 3778 1750 3779 1762
rect 3814 1734 3815 1758
rect 3817 1734 3819 1758
rect 3823 1734 3825 1758
rect 3827 1734 3828 1758
rect 3842 1728 3843 1752
rect 3845 1728 3847 1752
rect 3851 1728 3853 1752
rect 3855 1728 3856 1752
rect 3889 1735 3890 1759
rect 3892 1735 3900 1759
rect 3902 1735 3903 1759
rect 4091 1743 4092 1755
rect 4094 1743 4096 1755
rect 4100 1743 4102 1755
rect 4104 1743 4105 1755
rect 4125 1744 4126 1756
rect 4128 1744 4129 1756
rect 3775 1695 3776 1707
rect 3778 1695 3779 1707
rect 3939 1715 3940 1727
rect 3942 1715 3944 1727
rect 3948 1715 3950 1727
rect 3952 1715 3953 1727
rect 4071 1713 4072 1725
rect 4074 1713 4075 1725
rect 4105 1713 4106 1725
rect 4108 1713 4110 1725
rect 4114 1713 4116 1725
rect 4118 1713 4119 1725
rect 4160 1708 4161 1732
rect 4163 1708 4171 1732
rect 4173 1708 4174 1732
rect 4026 1669 4027 1693
rect 4029 1669 4037 1693
rect 4039 1669 4040 1693
rect 4194 1707 4195 1719
rect 4197 1707 4198 1719
rect 4238 1708 4239 1720
rect 4241 1708 4242 1720
rect 4277 1692 4278 1716
rect 4280 1692 4282 1716
rect 4286 1692 4288 1716
rect 4290 1692 4291 1716
rect 4305 1686 4306 1710
rect 4308 1686 4310 1710
rect 4314 1686 4316 1710
rect 4318 1686 4319 1710
rect 4392 1699 4407 1711
rect 4392 1690 4395 1699
rect 4403 1690 4407 1699
rect 4392 1687 4407 1690
rect 4409 1691 4427 1711
rect 4523 1701 4526 1710
rect 4534 1701 4538 1710
rect 4523 1698 4538 1701
rect 4540 1702 4558 1710
rect 4540 1698 4546 1702
rect 4555 1698 4558 1702
rect 4409 1687 4415 1691
rect 4424 1687 4427 1691
rect 4606 1690 4609 1699
rect 4617 1690 4621 1699
rect 4238 1653 4239 1665
rect 4241 1653 4242 1665
rect 3347 1623 3362 1635
rect 3347 1614 3350 1623
rect 3358 1614 3362 1623
rect 3347 1611 3362 1614
rect 3364 1615 3382 1635
rect 4606 1687 4621 1690
rect 4623 1691 4641 1699
rect 4623 1687 4629 1691
rect 4638 1687 4641 1691
rect 4685 1690 4686 1697
rect 4692 1690 4694 1697
rect 3478 1625 3481 1634
rect 3489 1625 3493 1634
rect 3478 1622 3493 1625
rect 3495 1626 3513 1634
rect 4412 1660 4427 1666
rect 4412 1651 4415 1660
rect 4424 1651 4427 1660
rect 4412 1644 4427 1651
rect 4429 1652 4447 1666
rect 4429 1648 4435 1652
rect 4444 1648 4447 1652
rect 4429 1644 4447 1648
rect 4685 1685 4694 1690
rect 4696 1690 4711 1697
rect 4696 1685 4699 1690
rect 4710 1685 4711 1690
rect 3495 1622 3501 1626
rect 3510 1622 3513 1626
rect 3364 1611 3370 1615
rect 3379 1611 3382 1615
rect 3561 1614 3564 1623
rect 3572 1614 3576 1623
rect 3561 1611 3576 1614
rect 3578 1615 3596 1623
rect 3578 1611 3584 1615
rect 3593 1611 3596 1615
rect 3640 1614 3641 1621
rect 3647 1614 3649 1621
rect 3367 1584 3382 1590
rect 3367 1575 3370 1584
rect 3379 1575 3382 1584
rect 3367 1568 3382 1575
rect 3384 1576 3402 1590
rect 3384 1572 3390 1576
rect 3399 1572 3402 1576
rect 3384 1568 3402 1572
rect 3640 1609 3649 1614
rect 3651 1614 3666 1621
rect 3651 1609 3654 1614
rect 3665 1609 3666 1614
rect 4026 1545 4027 1569
rect 4029 1545 4037 1569
rect 4039 1545 4040 1569
rect 3775 1531 3776 1543
rect 3778 1531 3779 1543
rect 3814 1515 3815 1539
rect 3817 1515 3819 1539
rect 3823 1515 3825 1539
rect 3827 1515 3828 1539
rect 3842 1509 3843 1533
rect 3845 1509 3847 1533
rect 3851 1509 3853 1533
rect 3855 1509 3856 1533
rect 3889 1516 3890 1540
rect 3892 1516 3900 1540
rect 3902 1516 3903 1540
rect 4087 1524 4088 1536
rect 4090 1524 4092 1536
rect 4096 1524 4098 1536
rect 4100 1524 4101 1536
rect 4121 1525 4122 1537
rect 4124 1525 4125 1537
rect 3337 1476 3352 1488
rect 3337 1467 3340 1476
rect 3348 1467 3352 1476
rect 3337 1464 3352 1467
rect 3354 1468 3372 1488
rect 3468 1478 3471 1487
rect 3479 1478 3483 1487
rect 3468 1475 3483 1478
rect 3485 1479 3503 1487
rect 3485 1475 3491 1479
rect 3500 1475 3503 1479
rect 3354 1464 3360 1468
rect 3369 1464 3372 1468
rect 3551 1467 3554 1476
rect 3562 1467 3566 1476
rect 3551 1464 3566 1467
rect 3568 1468 3586 1476
rect 3775 1476 3776 1488
rect 3778 1476 3779 1488
rect 3568 1464 3574 1468
rect 3583 1464 3586 1468
rect 3630 1467 3631 1474
rect 3637 1467 3639 1474
rect 3357 1437 3372 1443
rect 3357 1428 3360 1437
rect 3369 1428 3372 1437
rect 3357 1421 3372 1428
rect 3374 1429 3392 1443
rect 3374 1425 3380 1429
rect 3389 1425 3392 1429
rect 3374 1421 3392 1425
rect 3630 1462 3639 1467
rect 3641 1467 3656 1474
rect 3641 1462 3644 1467
rect 3655 1462 3656 1467
rect 3939 1496 3940 1508
rect 3942 1496 3944 1508
rect 3948 1496 3950 1508
rect 3952 1496 3953 1508
rect 4071 1494 4072 1506
rect 4074 1494 4075 1506
rect 4105 1494 4106 1506
rect 4108 1494 4110 1506
rect 4114 1494 4116 1506
rect 4118 1494 4119 1506
rect 4159 1489 4160 1513
rect 4162 1489 4170 1513
rect 4172 1489 4173 1513
rect 4026 1450 4027 1474
rect 4029 1450 4037 1474
rect 4039 1450 4040 1474
rect 4193 1488 4194 1500
rect 4196 1488 4197 1500
rect 4235 1489 4236 1501
rect 4238 1489 4239 1501
rect 4274 1473 4275 1497
rect 4277 1473 4279 1497
rect 4283 1473 4285 1497
rect 4287 1473 4288 1497
rect 4302 1467 4303 1491
rect 4305 1467 4307 1491
rect 4311 1467 4313 1491
rect 4315 1467 4316 1491
rect 4392 1486 4407 1498
rect 4392 1477 4395 1486
rect 4403 1477 4407 1486
rect 4392 1474 4407 1477
rect 4409 1478 4427 1498
rect 4523 1488 4526 1497
rect 4534 1488 4538 1497
rect 4523 1485 4538 1488
rect 4540 1489 4558 1497
rect 4540 1485 4546 1489
rect 4555 1485 4558 1489
rect 4409 1474 4415 1478
rect 4424 1474 4427 1478
rect 4606 1477 4609 1486
rect 4617 1477 4621 1486
rect 4235 1434 4236 1446
rect 4238 1434 4239 1446
rect 4606 1474 4621 1477
rect 4623 1478 4641 1486
rect 4623 1474 4629 1478
rect 4638 1474 4641 1478
rect 4685 1477 4686 1484
rect 4692 1477 4694 1484
rect 4412 1447 4427 1453
rect 4412 1438 4415 1447
rect 4424 1438 4427 1447
rect 4412 1431 4427 1438
rect 4429 1439 4447 1453
rect 4429 1435 4435 1439
rect 4444 1435 4447 1439
rect 4429 1431 4447 1435
rect 4685 1472 4694 1477
rect 4696 1477 4711 1484
rect 4696 1472 4699 1477
rect 4710 1472 4711 1477
rect 3338 1329 3353 1341
rect 3338 1320 3341 1329
rect 3349 1320 3353 1329
rect 3338 1317 3353 1320
rect 3355 1321 3373 1341
rect 3469 1331 3472 1340
rect 3480 1331 3484 1340
rect 3469 1328 3484 1331
rect 3486 1332 3504 1340
rect 3486 1328 3492 1332
rect 3501 1328 3504 1332
rect 3355 1317 3361 1321
rect 3370 1317 3373 1321
rect 3552 1320 3555 1329
rect 3563 1320 3567 1329
rect 3552 1317 3567 1320
rect 3569 1321 3587 1329
rect 3569 1317 3575 1321
rect 3584 1317 3587 1321
rect 3631 1320 3632 1327
rect 3638 1320 3640 1327
rect 3358 1290 3373 1296
rect 3358 1281 3361 1290
rect 3370 1281 3373 1290
rect 3358 1274 3373 1281
rect 3375 1282 3393 1296
rect 3375 1278 3381 1282
rect 3390 1278 3393 1282
rect 3375 1274 3393 1278
rect 3631 1315 3640 1320
rect 3642 1320 3657 1327
rect 4023 1322 4024 1346
rect 4026 1322 4034 1346
rect 4036 1322 4037 1346
rect 3642 1315 3645 1320
rect 3656 1315 3657 1320
rect 3775 1308 3776 1320
rect 3778 1308 3779 1320
rect 3814 1292 3815 1316
rect 3817 1292 3819 1316
rect 3823 1292 3825 1316
rect 3827 1292 3828 1316
rect 3842 1286 3843 1310
rect 3845 1286 3847 1310
rect 3851 1286 3853 1310
rect 3855 1286 3856 1310
rect 3889 1293 3890 1317
rect 3892 1293 3900 1317
rect 3902 1293 3903 1317
rect 4085 1301 4086 1313
rect 4088 1301 4090 1313
rect 4094 1301 4096 1313
rect 4098 1301 4099 1313
rect 4119 1302 4120 1314
rect 4122 1302 4123 1314
rect 4163 1305 4164 1317
rect 4166 1305 4168 1317
rect 4172 1305 4174 1317
rect 4176 1305 4177 1317
rect 4197 1306 4198 1318
rect 4200 1306 4201 1318
rect 4230 1306 4231 1318
rect 4233 1306 4235 1318
rect 4239 1306 4241 1318
rect 4243 1306 4244 1318
rect 4264 1307 4265 1319
rect 4267 1307 4268 1319
rect 4389 1296 4404 1308
rect 3775 1253 3776 1265
rect 3778 1253 3779 1265
rect 4389 1287 4392 1296
rect 4400 1287 4404 1296
rect 3939 1273 3940 1285
rect 3942 1273 3944 1285
rect 3948 1273 3950 1285
rect 3952 1273 3953 1285
rect 4068 1271 4069 1283
rect 4071 1271 4072 1283
rect 4102 1271 4103 1283
rect 4105 1271 4107 1283
rect 4111 1271 4113 1283
rect 4115 1271 4116 1283
rect 4150 1263 4151 1287
rect 4153 1263 4161 1287
rect 4163 1263 4164 1287
rect 4389 1284 4404 1287
rect 4406 1288 4424 1308
rect 4520 1298 4523 1307
rect 4531 1298 4535 1307
rect 4520 1295 4535 1298
rect 4537 1299 4555 1307
rect 4537 1295 4543 1299
rect 4552 1295 4555 1299
rect 4406 1284 4412 1288
rect 4421 1284 4424 1288
rect 4603 1287 4606 1296
rect 4614 1287 4618 1296
rect 4023 1227 4024 1251
rect 4026 1227 4034 1251
rect 4036 1227 4037 1251
rect 4184 1262 4185 1274
rect 4187 1262 4188 1274
rect 4217 1250 4218 1274
rect 4220 1250 4228 1274
rect 4230 1250 4231 1274
rect 4603 1284 4618 1287
rect 4620 1288 4638 1296
rect 4620 1284 4626 1288
rect 4635 1284 4638 1288
rect 4682 1287 4683 1294
rect 4689 1287 4691 1294
rect 4251 1249 4252 1261
rect 4254 1249 4255 1261
rect 4409 1257 4424 1263
rect 4409 1248 4412 1257
rect 4421 1248 4424 1257
rect 4409 1241 4424 1248
rect 4426 1249 4444 1263
rect 4426 1245 4432 1249
rect 4441 1245 4444 1249
rect 4426 1241 4444 1245
rect 4682 1282 4691 1287
rect 4693 1287 4708 1294
rect 4693 1282 4696 1287
rect 4707 1282 4708 1287
rect 3347 1167 3362 1179
rect 3347 1158 3350 1167
rect 3358 1158 3362 1167
rect 3347 1155 3362 1158
rect 3364 1159 3382 1179
rect 3478 1169 3481 1178
rect 3489 1169 3493 1178
rect 3478 1166 3493 1169
rect 3495 1170 3513 1178
rect 3495 1166 3501 1170
rect 3510 1166 3513 1170
rect 3364 1155 3370 1159
rect 3379 1155 3382 1159
rect 3561 1158 3564 1167
rect 3572 1158 3576 1167
rect 3561 1155 3576 1158
rect 3578 1159 3596 1167
rect 3578 1155 3584 1159
rect 3593 1155 3596 1159
rect 3640 1158 3641 1165
rect 3647 1158 3649 1165
rect 3367 1128 3382 1134
rect 3367 1119 3370 1128
rect 3379 1119 3382 1128
rect 3367 1112 3382 1119
rect 3384 1120 3402 1134
rect 3384 1116 3390 1120
rect 3399 1116 3402 1120
rect 3384 1112 3402 1116
rect 3640 1153 3649 1158
rect 3651 1158 3666 1165
rect 3651 1153 3654 1158
rect 3665 1153 3666 1158
rect 3349 1029 3364 1041
rect 3349 1020 3352 1029
rect 3360 1020 3364 1029
rect 3349 1017 3364 1020
rect 3366 1021 3384 1041
rect 3480 1031 3483 1040
rect 3491 1031 3495 1040
rect 3480 1028 3495 1031
rect 3497 1032 3515 1040
rect 3497 1028 3503 1032
rect 3512 1028 3515 1032
rect 3366 1017 3372 1021
rect 3381 1017 3384 1021
rect 3563 1020 3566 1029
rect 3574 1020 3578 1029
rect 3563 1017 3578 1020
rect 3580 1021 3598 1029
rect 3580 1017 3586 1021
rect 3595 1017 3598 1021
rect 3642 1020 3643 1027
rect 3649 1020 3651 1027
rect 3369 990 3384 996
rect 3369 981 3372 990
rect 3381 981 3384 990
rect 3369 974 3384 981
rect 3386 982 3404 996
rect 3386 978 3392 982
rect 3401 978 3404 982
rect 3386 974 3404 978
rect 3642 1015 3651 1020
rect 3653 1020 3668 1027
rect 3653 1015 3656 1020
rect 3667 1015 3668 1020
<< ndcontact >>
rect 4135 2154 4139 2160
rect 4143 2154 4147 2160
rect 4174 2142 4178 2154
rect 4192 2142 4196 2154
rect 4202 2142 4206 2154
rect 4220 2142 4224 2154
rect 4135 2099 4139 2105
rect 4143 2099 4147 2105
rect 4480 2107 4489 2112
rect 4500 2113 4509 2119
rect 4561 2107 4570 2112
rect 4583 2113 4592 2119
rect 4639 2087 4646 2091
rect 4653 2087 4664 2093
rect 4369 2070 4377 2075
rect 4389 2070 4398 2076
rect 4460 2075 4468 2080
rect 4480 2081 4489 2087
rect 4543 2075 4551 2080
rect 4561 2081 4570 2087
rect 3467 2038 3476 2043
rect 3487 2044 3496 2050
rect 3548 2038 3557 2043
rect 3570 2044 3579 2050
rect 3626 2018 3633 2022
rect 3640 2018 3651 2024
rect 3356 2001 3364 2006
rect 3376 2001 3385 2007
rect 3447 2006 3455 2011
rect 3467 2012 3476 2018
rect 3530 2006 3538 2011
rect 3548 2012 3557 2018
rect 3771 1971 3775 1977
rect 3779 1971 3783 1977
rect 4061 1966 4065 1972
rect 4069 1966 4073 1972
rect 4162 1980 4166 1986
rect 4170 1980 4174 1986
rect 4201 1968 4205 1980
rect 4219 1968 4223 1980
rect 4229 1968 4233 1980
rect 4247 1968 4251 1980
rect 4027 1960 4031 1966
rect 4036 1960 4040 1966
rect 4045 1960 4049 1966
rect 3885 1949 3889 1955
rect 3894 1949 3898 1955
rect 3903 1949 3907 1955
rect 4085 1954 4089 1966
rect 4103 1954 4107 1966
rect 3810 1922 3814 1934
rect 3828 1922 3832 1934
rect 3838 1922 3842 1934
rect 3856 1922 3860 1934
rect 3935 1924 3939 1936
rect 3953 1924 3957 1936
rect 4162 1925 4166 1931
rect 4170 1925 4174 1931
rect 3771 1916 3775 1922
rect 3779 1916 3783 1922
rect 3474 1885 3483 1890
rect 3494 1891 3503 1897
rect 3555 1885 3564 1890
rect 3577 1891 3586 1897
rect 4516 1908 4525 1913
rect 4536 1914 4545 1920
rect 4597 1908 4606 1913
rect 4619 1914 4628 1920
rect 4675 1888 4682 1892
rect 4689 1888 4700 1894
rect 4405 1871 4413 1876
rect 4425 1871 4434 1877
rect 4496 1876 4504 1881
rect 4516 1882 4525 1888
rect 4579 1876 4587 1881
rect 4597 1882 4606 1888
rect 3633 1865 3640 1869
rect 3647 1865 3658 1871
rect 3363 1848 3371 1853
rect 3383 1848 3392 1854
rect 3454 1853 3462 1858
rect 3474 1859 3483 1865
rect 3537 1853 3545 1858
rect 3555 1859 3564 1865
rect 3475 1734 3484 1739
rect 3495 1740 3504 1746
rect 3556 1734 3565 1739
rect 3578 1740 3587 1746
rect 4087 1775 4091 1787
rect 4105 1775 4109 1787
rect 3771 1730 3775 1736
rect 3779 1730 3783 1736
rect 4121 1770 4125 1776
rect 4129 1770 4133 1776
rect 4022 1737 4026 1743
rect 4031 1737 4035 1743
rect 4040 1737 4044 1743
rect 3634 1714 3641 1718
rect 3648 1714 3659 1720
rect 3364 1697 3372 1702
rect 3384 1697 3393 1703
rect 3455 1702 3463 1707
rect 3475 1708 3484 1714
rect 3538 1702 3546 1707
rect 3556 1708 3565 1714
rect 3885 1708 3889 1714
rect 3894 1708 3898 1714
rect 3903 1708 3907 1714
rect 4022 1714 4026 1720
rect 4031 1714 4035 1720
rect 4040 1714 4044 1720
rect 3810 1681 3814 1693
rect 3828 1681 3832 1693
rect 3838 1681 3842 1693
rect 3856 1681 3860 1693
rect 3935 1683 3939 1695
rect 3953 1683 3957 1695
rect 4067 1693 4071 1699
rect 4075 1693 4079 1699
rect 3771 1675 3775 1681
rect 3779 1675 3783 1681
rect 4101 1681 4105 1693
rect 4119 1681 4123 1693
rect 4190 1687 4194 1693
rect 4198 1687 4202 1693
rect 4234 1688 4238 1694
rect 4242 1688 4246 1694
rect 4156 1681 4160 1687
rect 4165 1681 4169 1687
rect 4174 1681 4178 1687
rect 4273 1639 4277 1651
rect 4291 1639 4295 1651
rect 4301 1639 4305 1651
rect 4319 1639 4323 1651
rect 4234 1633 4238 1639
rect 4242 1633 4246 1639
rect 4526 1655 4535 1660
rect 4546 1661 4555 1667
rect 4607 1655 4616 1660
rect 4629 1661 4638 1667
rect 4685 1635 4692 1639
rect 4699 1635 4710 1641
rect 4415 1618 4423 1623
rect 4435 1618 4444 1624
rect 4506 1623 4514 1628
rect 4526 1629 4535 1635
rect 4589 1623 4597 1628
rect 4607 1629 4616 1635
rect 3481 1579 3490 1584
rect 3501 1585 3510 1591
rect 3562 1579 3571 1584
rect 3584 1585 3593 1591
rect 3640 1559 3647 1563
rect 3654 1559 3665 1565
rect 3370 1542 3378 1547
rect 3390 1542 3399 1548
rect 3461 1547 3469 1552
rect 3481 1553 3490 1559
rect 3544 1547 3552 1552
rect 3562 1553 3571 1559
rect 4083 1556 4087 1568
rect 4101 1556 4105 1568
rect 3771 1511 3775 1517
rect 3779 1511 3783 1517
rect 4117 1551 4121 1557
rect 4125 1551 4129 1557
rect 4022 1518 4026 1524
rect 4031 1518 4035 1524
rect 4040 1518 4044 1524
rect 3885 1489 3889 1495
rect 3894 1489 3898 1495
rect 3903 1489 3907 1495
rect 4022 1495 4026 1501
rect 4031 1495 4035 1501
rect 4040 1495 4044 1501
rect 3810 1462 3814 1474
rect 3828 1462 3832 1474
rect 3838 1462 3842 1474
rect 3856 1462 3860 1474
rect 3935 1464 3939 1476
rect 3953 1464 3957 1476
rect 4067 1474 4071 1480
rect 4075 1474 4079 1480
rect 3471 1432 3480 1437
rect 3491 1438 3500 1444
rect 3552 1432 3561 1437
rect 3574 1438 3583 1444
rect 3771 1456 3775 1462
rect 3779 1456 3783 1462
rect 4101 1462 4105 1474
rect 4119 1462 4123 1474
rect 4189 1468 4193 1474
rect 4197 1468 4201 1474
rect 4231 1469 4235 1475
rect 4239 1469 4243 1475
rect 4155 1462 4159 1468
rect 4164 1462 4168 1468
rect 4173 1462 4177 1468
rect 4270 1420 4274 1432
rect 4288 1420 4292 1432
rect 4298 1420 4302 1432
rect 4316 1420 4320 1432
rect 3630 1412 3637 1416
rect 3644 1412 3655 1418
rect 4231 1414 4235 1420
rect 4239 1414 4243 1420
rect 4526 1442 4535 1447
rect 4546 1448 4555 1454
rect 4607 1442 4616 1447
rect 4629 1448 4638 1454
rect 4685 1422 4692 1426
rect 4699 1422 4710 1428
rect 3360 1395 3368 1400
rect 3380 1395 3389 1401
rect 3451 1400 3459 1405
rect 3471 1406 3480 1412
rect 3534 1400 3542 1405
rect 3552 1406 3561 1412
rect 4415 1405 4423 1410
rect 4435 1405 4444 1411
rect 4506 1410 4514 1415
rect 4526 1416 4535 1422
rect 4589 1410 4597 1415
rect 4607 1416 4616 1422
rect 4081 1333 4085 1345
rect 4099 1333 4103 1345
rect 4159 1337 4163 1349
rect 4177 1337 4181 1349
rect 4226 1338 4230 1350
rect 4244 1338 4248 1350
rect 3472 1285 3481 1290
rect 3492 1291 3501 1297
rect 3553 1285 3562 1290
rect 3575 1291 3584 1297
rect 3771 1288 3775 1294
rect 3779 1288 3783 1294
rect 4115 1328 4119 1334
rect 4123 1328 4127 1334
rect 4193 1332 4197 1338
rect 4201 1332 4205 1338
rect 4260 1333 4264 1339
rect 4268 1333 4272 1339
rect 4019 1295 4023 1301
rect 4028 1295 4032 1301
rect 4037 1295 4041 1301
rect 3631 1265 3638 1269
rect 3645 1265 3656 1271
rect 3361 1248 3369 1253
rect 3381 1248 3390 1254
rect 3452 1253 3460 1258
rect 3472 1259 3481 1265
rect 3535 1253 3543 1258
rect 3553 1259 3562 1265
rect 3885 1266 3889 1272
rect 3894 1266 3898 1272
rect 3903 1266 3907 1272
rect 4019 1272 4023 1278
rect 4028 1272 4032 1278
rect 4037 1272 4041 1278
rect 3810 1239 3814 1251
rect 3828 1239 3832 1251
rect 3838 1239 3842 1251
rect 3856 1239 3860 1251
rect 3935 1241 3939 1253
rect 3953 1241 3957 1253
rect 4064 1251 4068 1257
rect 4072 1251 4076 1257
rect 3771 1233 3775 1239
rect 3779 1233 3783 1239
rect 4098 1239 4102 1251
rect 4116 1239 4120 1251
rect 4180 1242 4184 1248
rect 4188 1242 4192 1248
rect 4146 1236 4150 1242
rect 4155 1236 4159 1242
rect 4164 1236 4168 1242
rect 4247 1229 4251 1235
rect 4255 1229 4259 1235
rect 4213 1223 4217 1229
rect 4222 1223 4226 1229
rect 4231 1223 4235 1229
rect 4523 1252 4532 1257
rect 4543 1258 4552 1264
rect 4604 1252 4613 1257
rect 4626 1258 4635 1264
rect 4682 1232 4689 1236
rect 4696 1232 4707 1238
rect 4412 1215 4420 1220
rect 4432 1215 4441 1221
rect 4503 1220 4511 1225
rect 4523 1226 4532 1232
rect 4586 1220 4594 1225
rect 4604 1226 4613 1232
rect 3481 1123 3490 1128
rect 3501 1129 3510 1135
rect 3562 1123 3571 1128
rect 3584 1129 3593 1135
rect 3640 1103 3647 1107
rect 3654 1103 3665 1109
rect 3370 1086 3378 1091
rect 3390 1086 3399 1092
rect 3461 1091 3469 1096
rect 3481 1097 3490 1103
rect 3544 1091 3552 1096
rect 3562 1097 3571 1103
rect 3483 985 3492 990
rect 3503 991 3512 997
rect 3564 985 3573 990
rect 3586 991 3595 997
rect 3642 965 3649 969
rect 3656 965 3667 971
rect 3372 948 3380 953
rect 3392 948 3401 954
rect 3463 953 3471 958
rect 3483 959 3492 965
rect 3546 953 3554 958
rect 3564 959 3573 965
<< pdcontact >>
rect 4349 2142 4357 2151
rect 4135 2128 4139 2140
rect 4143 2128 4147 2140
rect 4480 2153 4488 2162
rect 4500 2150 4509 2154
rect 4369 2139 4378 2143
rect 4563 2142 4571 2151
rect 3336 2073 3344 2082
rect 4583 2139 4592 2143
rect 4640 2142 4646 2149
rect 3467 2084 3475 2093
rect 3487 2081 3496 2085
rect 3356 2070 3365 2074
rect 3550 2073 3558 2082
rect 3570 2070 3579 2074
rect 3627 2073 3633 2080
rect 3356 2034 3365 2043
rect 3376 2031 3385 2035
rect 4135 2073 4139 2085
rect 4143 2073 4147 2085
rect 4174 2077 4178 2101
rect 4183 2077 4187 2101
rect 4192 2077 4196 2101
rect 4202 2083 4206 2107
rect 4211 2083 4215 2107
rect 4220 2083 4224 2107
rect 4369 2103 4378 2112
rect 4389 2100 4398 2104
rect 4653 2137 4664 2142
rect 3640 2068 3651 2073
rect 3771 1991 3775 2003
rect 3779 1991 3783 2003
rect 3810 1975 3814 1999
rect 3819 1975 3823 1999
rect 3828 1975 3832 1999
rect 3838 1969 3842 1993
rect 3847 1969 3851 1993
rect 3856 1969 3860 1993
rect 3885 1976 3889 2000
rect 3903 1976 3907 2000
rect 4027 1987 4031 2011
rect 4045 1987 4049 2011
rect 3343 1920 3351 1929
rect 3474 1931 3482 1940
rect 3771 1936 3775 1948
rect 3779 1936 3783 1948
rect 3494 1928 3503 1932
rect 3363 1917 3372 1921
rect 3557 1920 3565 1929
rect 3577 1917 3586 1921
rect 3634 1920 3640 1927
rect 3363 1881 3372 1890
rect 3383 1878 3392 1882
rect 3935 1956 3939 1968
rect 3944 1956 3948 1968
rect 3953 1956 3957 1968
rect 4061 1986 4065 1998
rect 4069 1986 4073 1998
rect 4085 1986 4089 1998
rect 4094 1986 4098 1998
rect 4103 1986 4107 1998
rect 4162 1954 4166 1966
rect 4170 1954 4174 1966
rect 4385 1943 4393 1952
rect 4516 1954 4524 1963
rect 4536 1951 4545 1955
rect 4405 1940 4414 1944
rect 4599 1943 4607 1952
rect 3647 1915 3658 1920
rect 4162 1899 4166 1911
rect 4170 1899 4174 1911
rect 4201 1903 4205 1927
rect 4210 1903 4214 1927
rect 4219 1903 4223 1927
rect 4229 1909 4233 1933
rect 4238 1909 4242 1933
rect 4247 1909 4251 1933
rect 4619 1940 4628 1944
rect 4676 1943 4682 1950
rect 4405 1904 4414 1913
rect 4425 1901 4434 1905
rect 4689 1938 4700 1943
rect 3344 1769 3352 1778
rect 3475 1780 3483 1789
rect 3495 1777 3504 1781
rect 3364 1766 3373 1770
rect 3558 1769 3566 1778
rect 3578 1766 3587 1770
rect 3635 1769 3641 1776
rect 3364 1730 3373 1739
rect 3384 1727 3393 1731
rect 3648 1764 3659 1769
rect 4022 1764 4026 1788
rect 4040 1764 4044 1788
rect 3771 1750 3775 1762
rect 3779 1750 3783 1762
rect 3810 1734 3814 1758
rect 3819 1734 3823 1758
rect 3828 1734 3832 1758
rect 3838 1728 3842 1752
rect 3847 1728 3851 1752
rect 3856 1728 3860 1752
rect 3885 1735 3889 1759
rect 3903 1735 3907 1759
rect 4087 1743 4091 1755
rect 4096 1743 4100 1755
rect 4105 1743 4109 1755
rect 4121 1744 4125 1756
rect 4129 1744 4133 1756
rect 3771 1695 3775 1707
rect 3779 1695 3783 1707
rect 3935 1715 3939 1727
rect 3944 1715 3948 1727
rect 3953 1715 3957 1727
rect 4067 1713 4071 1725
rect 4075 1713 4079 1725
rect 4101 1713 4105 1725
rect 4110 1713 4114 1725
rect 4119 1713 4123 1725
rect 4156 1708 4160 1732
rect 4174 1708 4178 1732
rect 4022 1669 4026 1693
rect 4040 1669 4044 1693
rect 4190 1707 4194 1719
rect 4198 1707 4202 1719
rect 4234 1708 4238 1720
rect 4242 1708 4246 1720
rect 4273 1692 4277 1716
rect 4282 1692 4286 1716
rect 4291 1692 4295 1716
rect 4301 1686 4305 1710
rect 4310 1686 4314 1710
rect 4319 1686 4323 1710
rect 4395 1690 4403 1699
rect 4526 1701 4534 1710
rect 4546 1698 4555 1702
rect 4415 1687 4424 1691
rect 4609 1690 4617 1699
rect 4234 1653 4238 1665
rect 4242 1653 4246 1665
rect 3350 1614 3358 1623
rect 4629 1687 4638 1691
rect 4686 1690 4692 1697
rect 3481 1625 3489 1634
rect 4415 1651 4424 1660
rect 4435 1648 4444 1652
rect 4699 1685 4710 1690
rect 3501 1622 3510 1626
rect 3370 1611 3379 1615
rect 3564 1614 3572 1623
rect 3584 1611 3593 1615
rect 3641 1614 3647 1621
rect 3370 1575 3379 1584
rect 3390 1572 3399 1576
rect 3654 1609 3665 1614
rect 4022 1545 4026 1569
rect 4040 1545 4044 1569
rect 3771 1531 3775 1543
rect 3779 1531 3783 1543
rect 3810 1515 3814 1539
rect 3819 1515 3823 1539
rect 3828 1515 3832 1539
rect 3838 1509 3842 1533
rect 3847 1509 3851 1533
rect 3856 1509 3860 1533
rect 3885 1516 3889 1540
rect 3903 1516 3907 1540
rect 4083 1524 4087 1536
rect 4092 1524 4096 1536
rect 4101 1524 4105 1536
rect 4117 1525 4121 1537
rect 4125 1525 4129 1537
rect 3340 1467 3348 1476
rect 3471 1478 3479 1487
rect 3491 1475 3500 1479
rect 3360 1464 3369 1468
rect 3554 1467 3562 1476
rect 3771 1476 3775 1488
rect 3779 1476 3783 1488
rect 3574 1464 3583 1468
rect 3631 1467 3637 1474
rect 3360 1428 3369 1437
rect 3380 1425 3389 1429
rect 3644 1462 3655 1467
rect 3935 1496 3939 1508
rect 3944 1496 3948 1508
rect 3953 1496 3957 1508
rect 4067 1494 4071 1506
rect 4075 1494 4079 1506
rect 4101 1494 4105 1506
rect 4110 1494 4114 1506
rect 4119 1494 4123 1506
rect 4155 1489 4159 1513
rect 4173 1489 4177 1513
rect 4022 1450 4026 1474
rect 4040 1450 4044 1474
rect 4189 1488 4193 1500
rect 4197 1488 4201 1500
rect 4231 1489 4235 1501
rect 4239 1489 4243 1501
rect 4270 1473 4274 1497
rect 4279 1473 4283 1497
rect 4288 1473 4292 1497
rect 4298 1467 4302 1491
rect 4307 1467 4311 1491
rect 4316 1467 4320 1491
rect 4395 1477 4403 1486
rect 4526 1488 4534 1497
rect 4546 1485 4555 1489
rect 4415 1474 4424 1478
rect 4609 1477 4617 1486
rect 4231 1434 4235 1446
rect 4239 1434 4243 1446
rect 4629 1474 4638 1478
rect 4686 1477 4692 1484
rect 4415 1438 4424 1447
rect 4435 1435 4444 1439
rect 4699 1472 4710 1477
rect 3341 1320 3349 1329
rect 3472 1331 3480 1340
rect 3492 1328 3501 1332
rect 3361 1317 3370 1321
rect 3555 1320 3563 1329
rect 3575 1317 3584 1321
rect 3632 1320 3638 1327
rect 3361 1281 3370 1290
rect 3381 1278 3390 1282
rect 4019 1322 4023 1346
rect 4037 1322 4041 1346
rect 3645 1315 3656 1320
rect 3771 1308 3775 1320
rect 3779 1308 3783 1320
rect 3810 1292 3814 1316
rect 3819 1292 3823 1316
rect 3828 1292 3832 1316
rect 3838 1286 3842 1310
rect 3847 1286 3851 1310
rect 3856 1286 3860 1310
rect 3885 1293 3889 1317
rect 3903 1293 3907 1317
rect 4081 1301 4085 1313
rect 4090 1301 4094 1313
rect 4099 1301 4103 1313
rect 4115 1302 4119 1314
rect 4123 1302 4127 1314
rect 4159 1305 4163 1317
rect 4168 1305 4172 1317
rect 4177 1305 4181 1317
rect 4193 1306 4197 1318
rect 4201 1306 4205 1318
rect 4226 1306 4230 1318
rect 4235 1306 4239 1318
rect 4244 1306 4248 1318
rect 4260 1307 4264 1319
rect 4268 1307 4272 1319
rect 3771 1253 3775 1265
rect 3779 1253 3783 1265
rect 4392 1287 4400 1296
rect 3935 1273 3939 1285
rect 3944 1273 3948 1285
rect 3953 1273 3957 1285
rect 4064 1271 4068 1283
rect 4072 1271 4076 1283
rect 4098 1271 4102 1283
rect 4107 1271 4111 1283
rect 4116 1271 4120 1283
rect 4146 1263 4150 1287
rect 4164 1263 4168 1287
rect 4523 1298 4531 1307
rect 4543 1295 4552 1299
rect 4412 1284 4421 1288
rect 4606 1287 4614 1296
rect 4019 1227 4023 1251
rect 4037 1227 4041 1251
rect 4180 1262 4184 1274
rect 4188 1262 4192 1274
rect 4213 1250 4217 1274
rect 4231 1250 4235 1274
rect 4626 1284 4635 1288
rect 4683 1287 4689 1294
rect 4247 1249 4251 1261
rect 4255 1249 4259 1261
rect 4412 1248 4421 1257
rect 4432 1245 4441 1249
rect 4696 1282 4707 1287
rect 3350 1158 3358 1167
rect 3481 1169 3489 1178
rect 3501 1166 3510 1170
rect 3370 1155 3379 1159
rect 3564 1158 3572 1167
rect 3584 1155 3593 1159
rect 3641 1158 3647 1165
rect 3370 1119 3379 1128
rect 3390 1116 3399 1120
rect 3654 1153 3665 1158
rect 3352 1020 3360 1029
rect 3483 1031 3491 1040
rect 3503 1028 3512 1032
rect 3372 1017 3381 1021
rect 3566 1020 3574 1029
rect 3586 1017 3595 1021
rect 3643 1020 3649 1027
rect 3372 981 3381 990
rect 3392 978 3401 982
rect 3656 1015 3667 1020
<< polysilicon >>
rect 4361 2163 4363 2175
rect 4140 2160 4142 2163
rect 4179 2154 4181 2157
rect 4189 2154 4191 2157
rect 4207 2154 4209 2157
rect 4217 2154 4219 2157
rect 4140 2140 4142 2154
rect 4140 2125 4142 2128
rect 4179 2115 4181 2142
rect 4189 2116 4191 2142
rect 4207 2122 4209 2142
rect 4217 2133 4219 2142
rect 4492 2162 4494 2170
rect 4575 2151 4577 2158
rect 4492 2142 4494 2150
rect 4459 2140 4494 2142
rect 3348 2094 3350 2106
rect 4140 2105 4142 2108
rect 3479 2093 3481 2101
rect 4179 2101 4181 2110
rect 4189 2101 4191 2111
rect 4207 2107 4209 2118
rect 4217 2107 4219 2129
rect 4361 2128 4363 2139
rect 4459 2131 4461 2140
rect 4648 2149 4650 2156
rect 4448 2129 4461 2131
rect 4346 2126 4363 2128
rect 3562 2082 3564 2089
rect 3479 2073 3481 2081
rect 3446 2071 3481 2073
rect 3348 2059 3350 2070
rect 3446 2062 3448 2071
rect 3635 2080 3637 2087
rect 4140 2085 4142 2099
rect 3435 2060 3448 2062
rect 3333 2057 3350 2059
rect 3333 2041 3335 2057
rect 3368 2049 3370 2060
rect 3321 2037 3335 2041
rect 3333 2016 3335 2037
rect 3333 2014 3353 2016
rect 3368 2014 3370 2027
rect 3435 2021 3437 2060
rect 3479 2050 3481 2064
rect 3562 2060 3564 2070
rect 4346 2110 4348 2126
rect 4381 2118 4383 2129
rect 4339 2106 4348 2110
rect 4346 2085 4348 2106
rect 4346 2083 4366 2085
rect 4381 2083 4383 2096
rect 4448 2090 4450 2129
rect 4492 2119 4494 2133
rect 4575 2129 4577 2139
rect 4547 2127 4577 2129
rect 4492 2101 4494 2107
rect 4547 2091 4549 2127
rect 4579 2119 4581 2122
rect 4579 2098 4581 2107
rect 4648 2093 4650 2137
rect 4448 2088 4474 2090
rect 4547 2089 4557 2091
rect 4472 2087 4474 2088
rect 4555 2087 4557 2089
rect 4207 2080 4209 2083
rect 4217 2080 4219 2083
rect 4364 2079 4366 2083
rect 4364 2077 4383 2079
rect 4179 2074 4181 2077
rect 4189 2074 4191 2077
rect 4381 2076 4383 2077
rect 4140 2070 4142 2073
rect 4648 2079 4650 2087
rect 3534 2058 3564 2060
rect 3479 2032 3481 2038
rect 3534 2022 3536 2058
rect 3566 2050 3568 2053
rect 3566 2029 3568 2038
rect 3635 2024 3637 2068
rect 4381 2064 4383 2070
rect 4472 2069 4474 2075
rect 4555 2069 4557 2075
rect 3435 2019 3461 2021
rect 3534 2020 3544 2022
rect 3459 2018 3461 2019
rect 3542 2018 3544 2020
rect 3351 2010 3353 2014
rect 3351 2008 3370 2010
rect 3368 2007 3370 2008
rect 3635 2010 3637 2018
rect 4032 2011 4034 2014
rect 4042 2011 4044 2014
rect 3368 1995 3370 2001
rect 3459 2000 3461 2006
rect 3542 2000 3544 2006
rect 3776 2003 3778 2006
rect 3815 1999 3817 2002
rect 3825 1999 3827 2002
rect 3890 2000 3892 2003
rect 3900 2000 3902 2003
rect 3776 1977 3778 1991
rect 3843 1993 3845 1996
rect 3853 1993 3855 1996
rect 3776 1968 3778 1971
rect 3815 1966 3817 1975
rect 3825 1965 3827 1975
rect 4066 1998 4068 2001
rect 4090 1998 4092 2001
rect 4100 1998 4102 2001
rect 3355 1941 3357 1953
rect 3776 1948 3778 1951
rect 3486 1940 3488 1948
rect 3569 1929 3571 1936
rect 3486 1920 3488 1928
rect 3453 1918 3488 1920
rect 3355 1906 3357 1917
rect 3453 1909 3455 1918
rect 3642 1927 3644 1934
rect 3442 1907 3455 1909
rect 3340 1904 3357 1906
rect 3340 1888 3342 1904
rect 3375 1896 3377 1907
rect 3328 1884 3342 1888
rect 3340 1863 3342 1884
rect 3340 1861 3360 1863
rect 3375 1861 3377 1874
rect 3442 1868 3444 1907
rect 3486 1897 3488 1911
rect 3569 1907 3571 1917
rect 3776 1922 3778 1936
rect 3815 1934 3817 1961
rect 3825 1934 3827 1960
rect 3843 1958 3845 1969
rect 3843 1934 3845 1954
rect 3853 1947 3855 1969
rect 3890 1955 3892 1976
rect 3900 1955 3902 1976
rect 3940 1968 3942 1971
rect 3950 1968 3952 1971
rect 4032 1966 4034 1987
rect 4042 1966 4044 1987
rect 4167 1986 4169 1989
rect 4066 1972 4068 1986
rect 4090 1966 4092 1986
rect 4100 1966 4102 1986
rect 4206 1980 4208 1983
rect 4216 1980 4218 1983
rect 4234 1980 4236 1983
rect 4244 1980 4246 1983
rect 4167 1966 4169 1980
rect 4066 1963 4068 1966
rect 4032 1957 4034 1960
rect 4042 1957 4044 1960
rect 3890 1946 3892 1949
rect 3900 1946 3902 1949
rect 3853 1934 3855 1943
rect 3940 1936 3942 1956
rect 3950 1936 3952 1956
rect 4090 1951 4092 1954
rect 4100 1951 4102 1954
rect 4167 1951 4169 1954
rect 4206 1941 4208 1968
rect 4216 1942 4218 1968
rect 4234 1948 4236 1968
rect 4244 1959 4246 1968
rect 4397 1964 4399 1976
rect 4167 1931 4169 1934
rect 4206 1927 4208 1936
rect 4216 1927 4218 1937
rect 4234 1933 4236 1944
rect 4244 1933 4246 1955
rect 4528 1963 4530 1971
rect 4611 1952 4613 1959
rect 4528 1943 4530 1951
rect 4495 1941 4530 1943
rect 3815 1919 3817 1922
rect 3825 1919 3827 1922
rect 3843 1919 3845 1922
rect 3853 1919 3855 1922
rect 3940 1921 3942 1924
rect 3950 1921 3952 1924
rect 3541 1905 3571 1907
rect 3486 1879 3488 1885
rect 3541 1869 3543 1905
rect 3573 1897 3575 1900
rect 3573 1876 3575 1885
rect 3642 1871 3644 1915
rect 3776 1913 3778 1916
rect 4167 1911 4169 1925
rect 4397 1929 4399 1940
rect 4495 1932 4497 1941
rect 4684 1950 4686 1957
rect 4484 1930 4497 1932
rect 4382 1927 4399 1929
rect 4382 1911 4384 1927
rect 4417 1919 4419 1930
rect 4234 1906 4236 1909
rect 4244 1906 4246 1909
rect 4378 1907 4384 1911
rect 4206 1900 4208 1903
rect 4216 1900 4218 1903
rect 4167 1896 4169 1899
rect 4382 1886 4384 1907
rect 4382 1884 4402 1886
rect 4417 1884 4419 1897
rect 4484 1891 4486 1930
rect 4528 1920 4530 1934
rect 4611 1930 4613 1940
rect 4583 1928 4613 1930
rect 4528 1902 4530 1908
rect 4583 1892 4585 1928
rect 4615 1920 4617 1923
rect 4615 1899 4617 1908
rect 4684 1894 4686 1938
rect 4484 1889 4510 1891
rect 4583 1890 4593 1892
rect 4508 1888 4510 1889
rect 4591 1888 4593 1890
rect 4400 1880 4402 1884
rect 4400 1878 4419 1880
rect 4417 1877 4419 1878
rect 4684 1880 4686 1888
rect 3442 1866 3468 1868
rect 3541 1867 3551 1869
rect 3466 1865 3468 1866
rect 3549 1865 3551 1867
rect 4417 1865 4419 1871
rect 4508 1870 4510 1876
rect 4591 1870 4593 1876
rect 3358 1857 3360 1861
rect 3358 1855 3377 1857
rect 3375 1854 3377 1855
rect 3642 1857 3644 1865
rect 3375 1842 3377 1848
rect 3466 1847 3468 1853
rect 3549 1847 3551 1853
rect 3356 1790 3358 1802
rect 3487 1789 3489 1797
rect 4027 1788 4029 1791
rect 4037 1788 4039 1791
rect 3570 1778 3572 1785
rect 3487 1769 3489 1777
rect 3454 1767 3489 1769
rect 3356 1755 3358 1766
rect 3454 1758 3456 1767
rect 3643 1776 3645 1783
rect 3443 1756 3456 1758
rect 3341 1753 3358 1755
rect 3341 1737 3343 1753
rect 3376 1745 3378 1756
rect 3329 1733 3343 1737
rect 3341 1712 3343 1733
rect 3341 1710 3361 1712
rect 3376 1710 3378 1723
rect 3443 1717 3445 1756
rect 3487 1746 3489 1760
rect 3570 1756 3572 1766
rect 3542 1754 3572 1756
rect 3487 1728 3489 1734
rect 3542 1718 3544 1754
rect 3574 1746 3576 1749
rect 3574 1725 3576 1734
rect 3643 1720 3645 1764
rect 3776 1762 3778 1765
rect 4092 1787 4094 1790
rect 4102 1787 4104 1790
rect 4126 1776 4128 1779
rect 3815 1758 3817 1761
rect 3825 1758 3827 1761
rect 3890 1759 3892 1762
rect 3900 1759 3902 1762
rect 3776 1736 3778 1750
rect 3843 1752 3845 1755
rect 3853 1752 3855 1755
rect 3776 1727 3778 1730
rect 3815 1725 3817 1734
rect 3825 1724 3827 1734
rect 4027 1743 4029 1764
rect 4037 1743 4039 1764
rect 4092 1755 4094 1775
rect 4102 1755 4104 1775
rect 4126 1756 4128 1770
rect 4092 1740 4094 1743
rect 4102 1740 4104 1743
rect 4126 1741 4128 1744
rect 3443 1715 3469 1717
rect 3542 1716 3552 1718
rect 3467 1714 3469 1715
rect 3550 1714 3552 1716
rect 3359 1706 3361 1710
rect 3359 1704 3378 1706
rect 3376 1703 3378 1704
rect 3643 1706 3645 1714
rect 3776 1707 3778 1710
rect 3376 1691 3378 1697
rect 3467 1696 3469 1702
rect 3550 1696 3552 1702
rect 3776 1681 3778 1695
rect 3815 1693 3817 1720
rect 3825 1693 3827 1719
rect 3843 1717 3845 1728
rect 3843 1693 3845 1713
rect 3853 1706 3855 1728
rect 3890 1714 3892 1735
rect 3900 1714 3902 1735
rect 4027 1734 4029 1737
rect 4037 1734 4039 1737
rect 4161 1732 4163 1735
rect 4171 1732 4173 1735
rect 3940 1727 3942 1730
rect 3950 1727 3952 1730
rect 4072 1725 4074 1728
rect 4106 1725 4108 1728
rect 4116 1725 4118 1728
rect 4027 1720 4029 1723
rect 4037 1720 4039 1723
rect 3890 1705 3892 1708
rect 3900 1705 3902 1708
rect 3853 1693 3855 1702
rect 3940 1695 3942 1715
rect 3950 1695 3952 1715
rect 4027 1693 4029 1714
rect 4037 1693 4039 1714
rect 4072 1699 4074 1713
rect 4106 1693 4108 1713
rect 4116 1693 4118 1713
rect 4195 1719 4197 1722
rect 4239 1720 4241 1723
rect 3815 1678 3817 1681
rect 3825 1678 3827 1681
rect 3843 1678 3845 1681
rect 3853 1678 3855 1681
rect 3940 1680 3942 1683
rect 3950 1680 3952 1683
rect 3776 1672 3778 1675
rect 4072 1690 4074 1693
rect 4161 1687 4163 1708
rect 4171 1687 4173 1708
rect 4278 1716 4280 1719
rect 4288 1716 4290 1719
rect 4195 1693 4197 1707
rect 4239 1694 4241 1708
rect 4306 1710 4308 1713
rect 4316 1710 4318 1713
rect 4407 1711 4409 1723
rect 4195 1684 4197 1687
rect 4239 1685 4241 1688
rect 4278 1683 4280 1692
rect 4106 1678 4108 1681
rect 4116 1678 4118 1681
rect 4161 1678 4163 1681
rect 4171 1678 4173 1681
rect 4288 1682 4290 1692
rect 4538 1710 4540 1718
rect 4621 1699 4623 1706
rect 4538 1690 4540 1698
rect 4505 1688 4540 1690
rect 4027 1666 4029 1669
rect 4037 1666 4039 1669
rect 4239 1665 4241 1668
rect 3362 1635 3364 1647
rect 3493 1634 3495 1642
rect 4239 1639 4241 1653
rect 4278 1651 4280 1678
rect 4288 1651 4290 1677
rect 4306 1675 4308 1686
rect 4306 1651 4308 1671
rect 4316 1664 4318 1686
rect 4407 1676 4409 1687
rect 4505 1679 4507 1688
rect 4694 1697 4696 1704
rect 4494 1677 4507 1679
rect 4392 1674 4409 1676
rect 4316 1651 4318 1660
rect 4392 1658 4394 1674
rect 4427 1666 4429 1677
rect 4386 1654 4394 1658
rect 4278 1636 4280 1639
rect 4288 1636 4290 1639
rect 4306 1636 4308 1639
rect 4316 1636 4318 1639
rect 4392 1633 4394 1654
rect 4239 1630 4241 1633
rect 4392 1631 4412 1633
rect 4427 1631 4429 1644
rect 4494 1638 4496 1677
rect 4538 1667 4540 1681
rect 4621 1677 4623 1687
rect 4593 1675 4623 1677
rect 4538 1649 4540 1655
rect 4593 1639 4595 1675
rect 4625 1667 4627 1670
rect 4625 1646 4627 1655
rect 4694 1641 4696 1685
rect 4494 1636 4520 1638
rect 4593 1637 4603 1639
rect 4518 1635 4520 1636
rect 4601 1635 4603 1637
rect 3576 1623 3578 1630
rect 3493 1614 3495 1622
rect 3460 1612 3495 1614
rect 3362 1600 3364 1611
rect 3460 1603 3462 1612
rect 3649 1621 3651 1628
rect 4410 1627 4412 1631
rect 4410 1625 4429 1627
rect 4427 1624 4429 1625
rect 3449 1601 3462 1603
rect 3347 1598 3364 1600
rect 3347 1582 3349 1598
rect 3382 1590 3384 1601
rect 3335 1578 3349 1582
rect 3347 1557 3349 1578
rect 3347 1555 3367 1557
rect 3382 1555 3384 1568
rect 3449 1562 3451 1601
rect 3493 1591 3495 1605
rect 3576 1601 3578 1611
rect 4694 1627 4696 1635
rect 4427 1612 4429 1618
rect 4518 1617 4520 1623
rect 4601 1617 4603 1623
rect 3548 1599 3578 1601
rect 3493 1573 3495 1579
rect 3548 1563 3550 1599
rect 3580 1591 3582 1594
rect 3580 1570 3582 1579
rect 3649 1565 3651 1609
rect 4027 1569 4029 1572
rect 4037 1569 4039 1572
rect 3449 1560 3475 1562
rect 3548 1561 3558 1563
rect 3473 1559 3475 1560
rect 3556 1559 3558 1561
rect 3365 1551 3367 1555
rect 3365 1549 3384 1551
rect 3382 1548 3384 1549
rect 3649 1551 3651 1559
rect 3382 1536 3384 1542
rect 3473 1541 3475 1547
rect 3556 1541 3558 1547
rect 3776 1543 3778 1546
rect 4088 1568 4090 1571
rect 4098 1568 4100 1571
rect 4122 1557 4124 1560
rect 3815 1539 3817 1542
rect 3825 1539 3827 1542
rect 3890 1540 3892 1543
rect 3900 1540 3902 1543
rect 3776 1517 3778 1531
rect 3843 1533 3845 1536
rect 3853 1533 3855 1536
rect 3776 1508 3778 1511
rect 3815 1506 3817 1515
rect 3825 1505 3827 1515
rect 4027 1524 4029 1545
rect 4037 1524 4039 1545
rect 4088 1536 4090 1556
rect 4098 1536 4100 1556
rect 4122 1537 4124 1551
rect 4088 1521 4090 1524
rect 4098 1521 4100 1524
rect 4122 1522 4124 1525
rect 3352 1488 3354 1500
rect 3483 1487 3485 1495
rect 3776 1488 3778 1491
rect 3566 1476 3568 1483
rect 3483 1467 3485 1475
rect 3450 1465 3485 1467
rect 3352 1453 3354 1464
rect 3450 1456 3452 1465
rect 3639 1474 3641 1481
rect 3439 1454 3452 1456
rect 3337 1451 3354 1453
rect 3337 1435 3339 1451
rect 3372 1443 3374 1454
rect 3325 1431 3339 1435
rect 3337 1410 3339 1431
rect 3337 1408 3357 1410
rect 3372 1408 3374 1421
rect 3439 1415 3441 1454
rect 3483 1444 3485 1458
rect 3566 1454 3568 1464
rect 3776 1462 3778 1476
rect 3815 1474 3817 1501
rect 3825 1474 3827 1500
rect 3843 1498 3845 1509
rect 3843 1474 3845 1494
rect 3853 1487 3855 1509
rect 3890 1495 3892 1516
rect 3900 1495 3902 1516
rect 4027 1515 4029 1518
rect 4037 1515 4039 1518
rect 4160 1513 4162 1516
rect 4170 1513 4172 1516
rect 3940 1508 3942 1511
rect 3950 1508 3952 1511
rect 4072 1506 4074 1509
rect 4106 1506 4108 1509
rect 4116 1506 4118 1509
rect 4027 1501 4029 1504
rect 4037 1501 4039 1504
rect 3890 1486 3892 1489
rect 3900 1486 3902 1489
rect 3853 1474 3855 1483
rect 3940 1476 3942 1496
rect 3950 1476 3952 1496
rect 4027 1474 4029 1495
rect 4037 1474 4039 1495
rect 4072 1480 4074 1494
rect 4106 1474 4108 1494
rect 4116 1474 4118 1494
rect 4194 1500 4196 1503
rect 4236 1501 4238 1504
rect 3538 1452 3568 1454
rect 3483 1426 3485 1432
rect 3538 1416 3540 1452
rect 3570 1444 3572 1447
rect 3570 1423 3572 1432
rect 3639 1418 3641 1462
rect 3815 1459 3817 1462
rect 3825 1459 3827 1462
rect 3843 1459 3845 1462
rect 3853 1459 3855 1462
rect 3940 1461 3942 1464
rect 3950 1461 3952 1464
rect 3776 1453 3778 1456
rect 4072 1471 4074 1474
rect 4160 1468 4162 1489
rect 4170 1468 4172 1489
rect 4275 1497 4277 1500
rect 4285 1497 4287 1500
rect 4407 1498 4409 1510
rect 4194 1474 4196 1488
rect 4236 1475 4238 1489
rect 4303 1491 4305 1494
rect 4313 1491 4315 1494
rect 4194 1465 4196 1468
rect 4236 1466 4238 1469
rect 4275 1464 4277 1473
rect 4106 1459 4108 1462
rect 4116 1459 4118 1462
rect 4160 1459 4162 1462
rect 4170 1459 4172 1462
rect 4285 1463 4287 1473
rect 4538 1497 4540 1505
rect 4621 1486 4623 1493
rect 4538 1477 4540 1485
rect 4505 1475 4540 1477
rect 4027 1447 4029 1450
rect 4037 1447 4039 1450
rect 4236 1446 4238 1449
rect 4236 1420 4238 1434
rect 4275 1432 4277 1459
rect 4285 1432 4287 1458
rect 4303 1456 4305 1467
rect 4303 1432 4305 1452
rect 4313 1445 4315 1467
rect 4407 1463 4409 1474
rect 4505 1466 4507 1475
rect 4694 1484 4696 1491
rect 4494 1464 4507 1466
rect 4392 1461 4409 1463
rect 4392 1445 4394 1461
rect 4427 1453 4429 1464
rect 4313 1432 4315 1441
rect 4388 1441 4394 1445
rect 4392 1420 4394 1441
rect 3439 1413 3465 1415
rect 3538 1414 3548 1416
rect 3463 1412 3465 1413
rect 3546 1412 3548 1414
rect 4275 1417 4277 1420
rect 4285 1417 4287 1420
rect 4303 1417 4305 1420
rect 4313 1417 4315 1420
rect 4392 1418 4412 1420
rect 4427 1418 4429 1431
rect 4494 1425 4496 1464
rect 4538 1454 4540 1468
rect 4621 1464 4623 1474
rect 4593 1462 4623 1464
rect 4538 1436 4540 1442
rect 4593 1426 4595 1462
rect 4625 1454 4627 1457
rect 4625 1433 4627 1442
rect 4694 1428 4696 1472
rect 4494 1423 4520 1425
rect 4593 1424 4603 1426
rect 4518 1422 4520 1423
rect 4601 1422 4603 1424
rect 4410 1414 4412 1418
rect 3355 1404 3357 1408
rect 3355 1402 3374 1404
rect 3372 1401 3374 1402
rect 3639 1404 3641 1412
rect 4236 1411 4238 1414
rect 4410 1412 4429 1414
rect 4427 1411 4429 1412
rect 4694 1414 4696 1422
rect 3372 1389 3374 1395
rect 3463 1394 3465 1400
rect 3546 1394 3548 1400
rect 4427 1399 4429 1405
rect 4518 1404 4520 1410
rect 4601 1404 4603 1410
rect 3353 1341 3355 1353
rect 4164 1349 4166 1352
rect 4174 1349 4176 1352
rect 4231 1350 4233 1353
rect 4241 1350 4243 1353
rect 3484 1340 3486 1348
rect 4024 1346 4026 1349
rect 4034 1346 4036 1349
rect 3567 1329 3569 1336
rect 3484 1320 3486 1328
rect 3451 1318 3486 1320
rect 3353 1306 3355 1317
rect 3451 1309 3453 1318
rect 3640 1327 3642 1334
rect 3440 1307 3453 1309
rect 3338 1304 3355 1306
rect 3338 1288 3340 1304
rect 3373 1296 3375 1307
rect 3326 1284 3340 1288
rect 3338 1263 3340 1284
rect 3338 1261 3358 1263
rect 3373 1261 3375 1274
rect 3440 1268 3442 1307
rect 3484 1297 3486 1311
rect 3567 1307 3569 1317
rect 3776 1320 3778 1323
rect 4086 1345 4088 1348
rect 4096 1345 4098 1348
rect 4198 1338 4200 1341
rect 4265 1339 4267 1342
rect 4120 1334 4122 1337
rect 3539 1305 3569 1307
rect 3484 1279 3486 1285
rect 3539 1269 3541 1305
rect 3571 1297 3573 1300
rect 3571 1276 3573 1285
rect 3640 1271 3642 1315
rect 3815 1316 3817 1319
rect 3825 1316 3827 1319
rect 3890 1317 3892 1320
rect 3900 1317 3902 1320
rect 3776 1294 3778 1308
rect 3843 1310 3845 1313
rect 3853 1310 3855 1313
rect 3776 1285 3778 1288
rect 3815 1283 3817 1292
rect 3825 1282 3827 1292
rect 4024 1301 4026 1322
rect 4034 1301 4036 1322
rect 4086 1313 4088 1333
rect 4096 1313 4098 1333
rect 4120 1314 4122 1328
rect 4164 1317 4166 1337
rect 4174 1317 4176 1337
rect 4198 1318 4200 1332
rect 4231 1318 4233 1338
rect 4241 1318 4243 1338
rect 4265 1319 4267 1333
rect 4404 1308 4406 1320
rect 4164 1302 4166 1305
rect 4174 1302 4176 1305
rect 4198 1303 4200 1306
rect 4231 1303 4233 1306
rect 4241 1303 4243 1306
rect 4265 1304 4267 1307
rect 4086 1298 4088 1301
rect 4096 1298 4098 1301
rect 4120 1299 4122 1302
rect 3440 1266 3466 1268
rect 3539 1267 3549 1269
rect 3464 1265 3466 1266
rect 3547 1265 3549 1267
rect 3776 1265 3778 1268
rect 3356 1257 3358 1261
rect 3356 1255 3375 1257
rect 3373 1254 3375 1255
rect 3640 1257 3642 1265
rect 3373 1242 3375 1248
rect 3464 1247 3466 1253
rect 3547 1247 3549 1253
rect 3776 1239 3778 1253
rect 3815 1251 3817 1278
rect 3825 1251 3827 1277
rect 3843 1275 3845 1286
rect 3843 1251 3845 1271
rect 3853 1264 3855 1286
rect 3890 1272 3892 1293
rect 3900 1272 3902 1293
rect 4024 1292 4026 1295
rect 4034 1292 4036 1295
rect 3940 1285 3942 1288
rect 3950 1285 3952 1288
rect 4151 1287 4153 1290
rect 4161 1287 4163 1290
rect 4069 1283 4071 1286
rect 4103 1283 4105 1286
rect 4113 1283 4115 1286
rect 4024 1278 4026 1281
rect 4034 1278 4036 1281
rect 3890 1263 3892 1266
rect 3900 1263 3902 1266
rect 3853 1251 3855 1260
rect 3940 1253 3942 1273
rect 3950 1253 3952 1273
rect 4024 1251 4026 1272
rect 4034 1251 4036 1272
rect 4069 1257 4071 1271
rect 4103 1251 4105 1271
rect 4113 1251 4115 1271
rect 4535 1307 4537 1315
rect 4618 1296 4620 1303
rect 4535 1287 4537 1295
rect 4502 1285 4537 1287
rect 4185 1274 4187 1277
rect 4218 1274 4220 1277
rect 4228 1274 4230 1277
rect 3815 1236 3817 1239
rect 3825 1236 3827 1239
rect 3843 1236 3845 1239
rect 3853 1236 3855 1239
rect 3940 1238 3942 1241
rect 3950 1238 3952 1241
rect 3776 1230 3778 1233
rect 4069 1248 4071 1251
rect 4151 1242 4153 1263
rect 4161 1242 4163 1263
rect 4185 1248 4187 1262
rect 4404 1273 4406 1284
rect 4502 1276 4504 1285
rect 4691 1294 4693 1301
rect 4491 1274 4504 1276
rect 4389 1271 4406 1273
rect 4252 1261 4254 1264
rect 4103 1236 4105 1239
rect 4113 1236 4115 1239
rect 4185 1239 4187 1242
rect 4151 1233 4153 1236
rect 4161 1233 4163 1236
rect 4218 1229 4220 1250
rect 4228 1229 4230 1250
rect 4389 1255 4391 1271
rect 4424 1263 4426 1274
rect 4384 1252 4391 1255
rect 4377 1251 4391 1252
rect 4252 1235 4254 1249
rect 4389 1230 4391 1251
rect 4024 1224 4026 1227
rect 4034 1224 4036 1227
rect 4252 1226 4254 1229
rect 4389 1228 4409 1230
rect 4424 1228 4426 1241
rect 4491 1235 4493 1274
rect 4535 1264 4537 1278
rect 4618 1274 4620 1284
rect 4590 1272 4620 1274
rect 4535 1246 4537 1252
rect 4590 1236 4592 1272
rect 4622 1264 4624 1267
rect 4622 1243 4624 1252
rect 4691 1238 4693 1282
rect 4491 1233 4517 1235
rect 4590 1234 4600 1236
rect 4515 1232 4517 1233
rect 4598 1232 4600 1234
rect 4407 1224 4409 1228
rect 4218 1220 4220 1223
rect 4228 1220 4230 1223
rect 4407 1222 4426 1224
rect 4424 1221 4426 1222
rect 4691 1224 4693 1232
rect 4424 1209 4426 1215
rect 4515 1214 4517 1220
rect 4598 1214 4600 1220
rect 3362 1179 3364 1191
rect 3493 1178 3495 1186
rect 3576 1167 3578 1174
rect 3493 1158 3495 1166
rect 3460 1156 3495 1158
rect 3362 1144 3364 1155
rect 3460 1147 3462 1156
rect 3649 1165 3651 1172
rect 3449 1145 3462 1147
rect 3347 1142 3364 1144
rect 3347 1126 3349 1142
rect 3382 1134 3384 1145
rect 3335 1122 3349 1126
rect 3347 1101 3349 1122
rect 3347 1099 3367 1101
rect 3382 1099 3384 1112
rect 3449 1106 3451 1145
rect 3493 1135 3495 1149
rect 3576 1145 3578 1155
rect 3548 1143 3578 1145
rect 3493 1117 3495 1123
rect 3548 1107 3550 1143
rect 3580 1135 3582 1138
rect 3580 1114 3582 1123
rect 3649 1109 3651 1153
rect 3449 1104 3475 1106
rect 3548 1105 3558 1107
rect 3473 1103 3475 1104
rect 3556 1103 3558 1105
rect 3365 1095 3367 1099
rect 3365 1093 3384 1095
rect 3382 1092 3384 1093
rect 3649 1095 3651 1103
rect 3382 1080 3384 1086
rect 3473 1085 3475 1091
rect 3556 1085 3558 1091
rect 3364 1041 3366 1053
rect 3495 1040 3497 1048
rect 3578 1029 3580 1036
rect 3495 1020 3497 1028
rect 3462 1018 3497 1020
rect 3364 1006 3366 1017
rect 3462 1009 3464 1018
rect 3651 1027 3653 1034
rect 3451 1007 3464 1009
rect 3349 1004 3366 1006
rect 3349 988 3351 1004
rect 3384 996 3386 1007
rect 3337 984 3351 988
rect 3349 963 3351 984
rect 3349 961 3369 963
rect 3384 961 3386 974
rect 3451 968 3453 1007
rect 3495 997 3497 1011
rect 3578 1007 3580 1017
rect 3550 1005 3580 1007
rect 3495 979 3497 985
rect 3550 969 3552 1005
rect 3582 997 3584 1000
rect 3582 976 3584 985
rect 3651 971 3653 1015
rect 3451 966 3477 968
rect 3550 967 3560 969
rect 3475 965 3477 966
rect 3558 965 3560 967
rect 3367 957 3369 961
rect 3367 955 3386 957
rect 3384 954 3386 955
rect 3651 957 3653 965
rect 3384 942 3386 948
rect 3475 947 3477 953
rect 3558 947 3560 953
<< polycontact >>
rect 4136 2147 4140 2151
rect 4216 2129 4220 2133
rect 4205 2118 4209 2122
rect 4136 2092 4140 2096
rect 3364 2014 3368 2018
rect 3475 2051 3479 2055
rect 4334 2105 4339 2111
rect 4377 2083 4381 2087
rect 4488 2120 4492 2124
rect 4542 2122 4547 2127
rect 4575 2098 4579 2102
rect 4644 2105 4648 2110
rect 4450 2084 4454 2088
rect 3529 2053 3534 2058
rect 3562 2029 3566 2033
rect 3631 2036 3635 2041
rect 3437 2015 3441 2019
rect 3772 1980 3776 1984
rect 3371 1861 3375 1865
rect 3482 1898 3486 1902
rect 3772 1925 3776 1929
rect 3841 1954 3845 1958
rect 3886 1958 3890 1962
rect 3896 1965 3900 1969
rect 4028 1969 4032 1973
rect 4038 1976 4042 1980
rect 4062 1975 4066 1979
rect 4086 1975 4090 1979
rect 4096 1969 4100 1973
rect 4163 1973 4167 1977
rect 3852 1943 3856 1947
rect 3936 1945 3940 1949
rect 3946 1939 3950 1943
rect 4243 1955 4247 1959
rect 4232 1944 4236 1948
rect 4163 1918 4167 1922
rect 3536 1900 3541 1905
rect 3569 1876 3573 1880
rect 3638 1883 3642 1888
rect 4370 1905 4378 1911
rect 4413 1884 4417 1888
rect 4524 1921 4528 1925
rect 4578 1923 4583 1928
rect 4611 1899 4615 1903
rect 4680 1906 4684 1911
rect 4486 1885 4490 1889
rect 3444 1862 3448 1866
rect 3372 1710 3376 1714
rect 3483 1747 3487 1751
rect 3537 1749 3542 1754
rect 3570 1725 3574 1729
rect 3639 1732 3643 1737
rect 3772 1739 3776 1743
rect 4023 1746 4027 1750
rect 4033 1753 4037 1757
rect 4088 1762 4092 1766
rect 4098 1768 4102 1772
rect 4122 1763 4126 1767
rect 3445 1711 3449 1715
rect 3772 1684 3776 1688
rect 3841 1713 3845 1717
rect 3886 1717 3890 1721
rect 3896 1724 3900 1728
rect 3852 1702 3856 1706
rect 3936 1704 3940 1708
rect 3946 1698 3950 1702
rect 4023 1707 4027 1711
rect 4033 1700 4037 1704
rect 4068 1702 4072 1706
rect 4102 1702 4106 1706
rect 4112 1696 4116 1700
rect 4157 1690 4161 1694
rect 4167 1697 4171 1701
rect 4191 1696 4195 1700
rect 4235 1697 4239 1701
rect 4235 1642 4239 1646
rect 4304 1671 4308 1675
rect 4315 1660 4319 1664
rect 4379 1654 4386 1658
rect 4423 1631 4427 1635
rect 4534 1668 4538 1672
rect 4588 1670 4593 1675
rect 4621 1646 4625 1650
rect 4690 1653 4694 1658
rect 4496 1632 4500 1636
rect 3378 1555 3382 1559
rect 3489 1592 3493 1596
rect 3543 1594 3548 1599
rect 3576 1570 3580 1574
rect 3645 1577 3649 1582
rect 3451 1556 3455 1560
rect 3772 1520 3776 1524
rect 4023 1527 4027 1531
rect 4033 1534 4037 1538
rect 4084 1543 4088 1547
rect 4094 1549 4098 1553
rect 4118 1544 4122 1548
rect 3368 1408 3372 1412
rect 3479 1445 3483 1449
rect 3772 1465 3776 1469
rect 3841 1494 3845 1498
rect 3886 1498 3890 1502
rect 3896 1505 3900 1509
rect 3852 1483 3856 1487
rect 3936 1485 3940 1489
rect 3946 1479 3950 1483
rect 4023 1488 4027 1492
rect 4033 1481 4037 1485
rect 4068 1483 4072 1487
rect 4102 1483 4106 1487
rect 4112 1477 4116 1481
rect 3533 1447 3538 1452
rect 3566 1423 3570 1427
rect 3635 1430 3639 1435
rect 4156 1471 4160 1475
rect 4166 1478 4170 1482
rect 4190 1477 4194 1481
rect 4232 1478 4236 1482
rect 4232 1423 4236 1427
rect 4301 1452 4305 1456
rect 4312 1441 4316 1445
rect 4379 1440 4388 1445
rect 3441 1409 3445 1413
rect 4423 1418 4427 1422
rect 4534 1455 4538 1459
rect 4588 1457 4593 1462
rect 4621 1433 4625 1437
rect 4690 1440 4694 1445
rect 4496 1419 4500 1423
rect 3369 1261 3373 1265
rect 3480 1298 3484 1302
rect 3534 1300 3539 1305
rect 3567 1276 3571 1280
rect 3636 1283 3640 1288
rect 3772 1297 3776 1301
rect 4020 1304 4024 1308
rect 4030 1311 4034 1315
rect 4082 1320 4086 1324
rect 4092 1326 4096 1330
rect 4116 1321 4120 1325
rect 4160 1324 4164 1328
rect 4170 1330 4174 1334
rect 4194 1325 4198 1329
rect 4227 1325 4231 1329
rect 4237 1331 4241 1335
rect 4261 1326 4265 1330
rect 3442 1262 3446 1266
rect 3772 1242 3776 1246
rect 3841 1271 3845 1275
rect 3886 1275 3890 1279
rect 3896 1282 3900 1286
rect 3852 1260 3856 1264
rect 3936 1262 3940 1266
rect 3946 1256 3950 1260
rect 4020 1265 4024 1269
rect 4030 1258 4034 1262
rect 4065 1260 4069 1264
rect 4099 1260 4103 1264
rect 4109 1254 4113 1258
rect 4147 1245 4151 1249
rect 4157 1252 4161 1256
rect 4181 1251 4185 1255
rect 4214 1232 4218 1236
rect 4224 1239 4228 1243
rect 4368 1252 4384 1259
rect 4248 1238 4252 1242
rect 4420 1228 4424 1232
rect 4531 1265 4535 1269
rect 4585 1267 4590 1272
rect 4618 1243 4622 1247
rect 4687 1250 4691 1255
rect 4493 1229 4497 1233
rect 3378 1099 3382 1103
rect 3489 1136 3493 1140
rect 3543 1138 3548 1143
rect 3576 1114 3580 1118
rect 3645 1121 3649 1126
rect 3451 1100 3455 1104
rect 3380 961 3384 965
rect 3491 998 3495 1002
rect 3545 1000 3550 1005
rect 3578 976 3582 980
rect 3647 983 3651 988
rect 3453 962 3457 966
<< metal1 >>
rect 3826 2199 3893 2202
rect 3898 2199 4025 2202
rect 4030 2199 4129 2202
rect 4134 2199 4229 2202
rect 3826 2175 4063 2178
rect 4339 2177 4405 2186
rect 4461 2179 4540 2180
rect 4060 2122 4063 2175
rect 4129 2164 4159 2167
rect 4135 2160 4138 2164
rect 4156 2161 4159 2164
rect 4156 2158 4161 2161
rect 4166 2158 4230 2161
rect 4103 2148 4121 2151
rect 4103 2124 4106 2148
rect 4144 2151 4147 2154
rect 4174 2154 4177 2158
rect 4221 2154 4224 2158
rect 4126 2148 4136 2151
rect 4144 2148 4159 2151
rect 4144 2140 4147 2148
rect 3826 2119 4012 2122
rect 3326 2108 3392 2117
rect 3448 2110 3527 2111
rect 3336 2082 3344 2108
rect 3384 2100 3392 2108
rect 3440 2102 3527 2110
rect 3440 2100 3448 2102
rect 3384 2091 3448 2100
rect 3467 2093 3475 2102
rect 3518 2100 3527 2102
rect 3518 2091 3677 2100
rect 3518 2090 3527 2091
rect 3356 2043 3365 2070
rect 3487 2058 3496 2081
rect 3550 2082 3558 2091
rect 3627 2080 3633 2091
rect 3570 2059 3579 2070
rect 3421 2051 3475 2055
rect 3487 2053 3529 2058
rect 3570 2053 3610 2059
rect 3376 2021 3385 2031
rect 3421 2021 3428 2051
rect 3487 2050 3496 2053
rect 3570 2050 3579 2053
rect 3361 2014 3364 2018
rect 3376 2016 3428 2021
rect 3376 2007 3385 2016
rect 3437 2011 3441 2015
rect 3467 2018 3476 2038
rect 3548 2018 3557 2038
rect 3605 2041 3610 2053
rect 3640 2044 3651 2068
rect 3605 2036 3631 2041
rect 3640 2035 3713 2044
rect 3560 2029 3562 2033
rect 3640 2024 3651 2035
rect 3701 2034 3713 2035
rect 3356 1988 3364 2001
rect 3447 1988 3455 2006
rect 3530 1988 3538 2006
rect 3626 1988 3633 2018
rect 3329 1978 3650 1988
rect 3702 1983 3713 2034
rect 3757 2018 3872 2020
rect 3757 2017 3926 2018
rect 3757 1983 3760 2017
rect 3869 2015 3926 2017
rect 3770 2009 3798 2012
rect 3771 2003 3774 2009
rect 3795 2008 3798 2009
rect 3795 2005 3853 2008
rect 3858 2005 3866 2008
rect 3702 1978 3757 1983
rect 3762 1980 3772 1983
rect 3780 1983 3783 1991
rect 3810 1999 3813 2005
rect 3829 1999 3832 2005
rect 3780 1980 3801 1983
rect 3780 1977 3783 1980
rect 3771 1967 3774 1971
rect 3765 1965 3789 1967
rect 3765 1964 3783 1965
rect 3333 1955 3399 1964
rect 3455 1957 3534 1958
rect 3343 1929 3351 1955
rect 3391 1947 3399 1955
rect 3447 1949 3534 1957
rect 3788 1964 3789 1965
rect 3798 1957 3801 1980
rect 3839 1999 3859 2002
rect 3839 1993 3842 1999
rect 3856 1993 3859 1999
rect 3820 1972 3823 1975
rect 3820 1969 3838 1972
rect 3848 1962 3851 1969
rect 3869 1968 3872 2015
rect 3879 2006 3893 2009
rect 3898 2006 3913 2009
rect 3885 2000 3888 2006
rect 3869 1965 3896 1968
rect 3904 1967 3907 1976
rect 3904 1964 3910 1967
rect 3848 1959 3865 1962
rect 3770 1956 3789 1957
rect 3765 1954 3789 1956
rect 3798 1954 3841 1957
rect 3447 1947 3455 1949
rect 3391 1938 3455 1947
rect 3474 1940 3482 1949
rect 3525 1947 3534 1949
rect 3771 1948 3774 1954
rect 3525 1938 3684 1947
rect 3525 1937 3534 1938
rect 3363 1890 3372 1917
rect 3494 1905 3503 1928
rect 3557 1929 3565 1938
rect 3634 1927 3640 1938
rect 3827 1943 3852 1946
rect 3827 1941 3830 1943
rect 3733 1925 3757 1928
rect 3577 1906 3586 1917
rect 3428 1898 3482 1902
rect 3494 1900 3536 1905
rect 3577 1900 3617 1906
rect 3383 1868 3392 1878
rect 3428 1868 3435 1898
rect 3494 1897 3503 1900
rect 3577 1897 3586 1900
rect 3368 1861 3371 1865
rect 3383 1863 3435 1868
rect 3383 1854 3392 1863
rect 3444 1858 3448 1862
rect 3474 1865 3483 1885
rect 3555 1865 3564 1885
rect 3612 1888 3617 1900
rect 3647 1891 3658 1915
rect 3733 1891 3742 1925
rect 3762 1925 3772 1928
rect 3780 1928 3783 1936
rect 3792 1938 3830 1941
rect 3862 1940 3865 1959
rect 3873 1959 3886 1962
rect 3792 1928 3795 1938
rect 3833 1937 3865 1940
rect 3833 1934 3836 1937
rect 3780 1925 3795 1928
rect 3759 1906 3762 1924
rect 3780 1922 3783 1925
rect 3832 1931 3838 1934
rect 3771 1912 3774 1916
rect 3792 1915 3797 1918
rect 3810 1918 3813 1922
rect 3857 1920 3860 1922
rect 3857 1918 3858 1920
rect 3802 1915 3858 1918
rect 3863 1915 3866 1918
rect 3792 1912 3795 1915
rect 3765 1909 3795 1912
rect 3873 1911 3876 1959
rect 3904 1961 3907 1964
rect 3895 1958 3907 1961
rect 3895 1955 3898 1958
rect 3885 1943 3888 1949
rect 3904 1943 3907 1949
rect 3923 1948 3926 2015
rect 3974 2000 3977 2093
rect 4009 2051 4012 2119
rect 4060 2119 4101 2122
rect 4156 2138 4159 2148
rect 4196 2142 4202 2145
rect 4349 2151 4357 2177
rect 4397 2169 4405 2177
rect 4453 2171 4540 2179
rect 4453 2169 4461 2171
rect 4397 2160 4461 2169
rect 4480 2162 4488 2171
rect 4531 2169 4540 2171
rect 4531 2160 4690 2169
rect 4531 2159 4540 2160
rect 4197 2139 4200 2142
rect 4156 2135 4194 2138
rect 4197 2136 4229 2139
rect 4191 2133 4194 2135
rect 4191 2130 4216 2133
rect 4226 2132 4229 2136
rect 4226 2129 4323 2132
rect 4226 2128 4230 2129
rect 4135 2122 4138 2128
rect 4129 2120 4153 2122
rect 4060 2113 4063 2119
rect 4134 2119 4153 2120
rect 4162 2119 4205 2122
rect 4129 2111 4147 2112
rect 4152 2111 4153 2112
rect 4129 2109 4153 2111
rect 4135 2105 4138 2109
rect 4033 2094 4121 2097
rect 4144 2096 4147 2099
rect 4162 2096 4165 2119
rect 4226 2117 4229 2128
rect 4212 2114 4229 2117
rect 4212 2107 4215 2114
rect 4311 2111 4323 2129
rect 4369 2112 4378 2139
rect 4500 2127 4509 2150
rect 4563 2151 4571 2160
rect 4640 2149 4646 2160
rect 4583 2128 4592 2139
rect 4311 2108 4334 2111
rect 4184 2104 4202 2107
rect 4184 2101 4187 2104
rect 4126 2093 4136 2096
rect 4144 2093 4165 2096
rect 4144 2085 4147 2093
rect 4312 2105 4334 2108
rect 4434 2120 4488 2124
rect 4500 2122 4542 2127
rect 4583 2122 4623 2128
rect 4389 2090 4398 2100
rect 4434 2090 4441 2120
rect 4500 2119 4509 2122
rect 4583 2119 4592 2122
rect 4374 2083 4377 2087
rect 4389 2085 4441 2090
rect 4135 2067 4138 2073
rect 4174 2071 4177 2077
rect 4193 2071 4196 2077
rect 4203 2077 4206 2083
rect 4220 2077 4223 2083
rect 4203 2074 4223 2077
rect 4389 2076 4398 2085
rect 4450 2080 4454 2084
rect 4480 2087 4489 2107
rect 4561 2087 4570 2107
rect 4618 2110 4623 2122
rect 4653 2113 4664 2137
rect 4618 2105 4644 2110
rect 4653 2105 4679 2113
rect 4573 2098 4575 2102
rect 4653 2093 4664 2105
rect 4159 2068 4230 2071
rect 4159 2067 4162 2068
rect 4134 2064 4162 2067
rect 4369 2057 4377 2070
rect 4460 2057 4468 2075
rect 4543 2057 4551 2075
rect 4639 2057 4646 2087
rect 4009 2048 4018 2051
rect 3971 1997 3977 2000
rect 4015 1979 4018 2048
rect 4342 2047 4663 2057
rect 4021 2017 4024 2020
rect 4029 2017 4060 2020
rect 4027 2011 4030 2017
rect 4057 2007 4060 2017
rect 4055 2004 4119 2007
rect 3929 1974 3963 1977
rect 4015 1976 4038 1979
rect 4046 1978 4049 1987
rect 4061 1998 4064 2004
rect 4085 1998 4088 2004
rect 4104 1998 4107 2004
rect 4154 1990 4186 1993
rect 4162 1986 4165 1990
rect 4183 1987 4186 1990
rect 4046 1975 4062 1978
rect 4070 1978 4073 1986
rect 4094 1983 4097 1986
rect 4094 1980 4107 1983
rect 4183 1984 4188 1987
rect 4193 1984 4257 1987
rect 4070 1975 4086 1978
rect 4104 1977 4107 1980
rect 3935 1968 3938 1974
rect 3954 1968 3957 1974
rect 3971 1970 4003 1973
rect 4008 1970 4028 1973
rect 4046 1972 4049 1975
rect 4070 1972 4073 1975
rect 4104 1974 4114 1977
rect 4037 1969 4049 1972
rect 4037 1966 4040 1969
rect 4082 1969 4096 1972
rect 4104 1966 4107 1974
rect 4119 1974 4148 1977
rect 4171 1977 4174 1980
rect 4201 1980 4204 1984
rect 4248 1980 4251 1984
rect 4153 1974 4163 1977
rect 4171 1974 4186 1977
rect 4171 1966 4174 1974
rect 4061 1962 4064 1966
rect 3944 1953 3947 1956
rect 4027 1954 4030 1960
rect 4046 1954 4049 1960
rect 4052 1959 4079 1962
rect 4052 1954 4055 1959
rect 3944 1950 3957 1953
rect 4021 1951 4055 1954
rect 3923 1945 3936 1948
rect 3954 1947 3957 1950
rect 3954 1944 3996 1947
rect 3879 1940 3916 1943
rect 3895 1934 3898 1940
rect 3919 1939 3946 1942
rect 3919 1911 3922 1939
rect 3954 1936 3957 1944
rect 4001 1944 4067 1947
rect 4076 1948 4079 1959
rect 4183 1964 4186 1974
rect 4223 1968 4229 1971
rect 4375 1978 4441 1987
rect 4497 1980 4576 1981
rect 4224 1965 4227 1968
rect 4183 1961 4221 1964
rect 4224 1962 4256 1965
rect 4218 1959 4221 1961
rect 4218 1956 4243 1959
rect 4253 1958 4256 1962
rect 4323 1958 4335 1959
rect 4253 1955 4335 1958
rect 4253 1954 4257 1955
rect 4085 1948 4088 1954
rect 4076 1945 4101 1948
rect 4106 1945 4122 1948
rect 4162 1948 4165 1954
rect 4156 1946 4180 1948
rect 4161 1945 4180 1946
rect 4189 1945 4232 1948
rect 4156 1937 4174 1938
rect 4179 1937 4180 1938
rect 4156 1935 4180 1937
rect 4162 1931 4165 1935
rect 3935 1920 3938 1924
rect 3929 1915 3931 1918
rect 3936 1918 3938 1920
rect 4136 1920 4148 1923
rect 3936 1915 3963 1918
rect 3798 1908 3922 1911
rect 3798 1906 3801 1908
rect 3759 1903 3801 1906
rect 3612 1883 3638 1888
rect 3647 1883 3742 1891
rect 3567 1876 3569 1880
rect 3647 1871 3658 1883
rect 3363 1835 3371 1848
rect 3454 1835 3462 1853
rect 3537 1835 3545 1853
rect 3633 1835 3640 1865
rect 4136 1859 4139 1920
rect 4171 1922 4174 1925
rect 4189 1922 4192 1945
rect 4253 1943 4256 1954
rect 4261 1952 4335 1955
rect 4239 1940 4256 1943
rect 4239 1933 4242 1940
rect 4211 1930 4229 1933
rect 4211 1927 4214 1930
rect 4153 1919 4163 1922
rect 4171 1919 4192 1922
rect 4171 1911 4174 1919
rect 4323 1912 4335 1952
rect 4385 1952 4393 1978
rect 4433 1970 4441 1978
rect 4489 1972 4576 1980
rect 4489 1970 4497 1972
rect 4433 1961 4497 1970
rect 4516 1963 4524 1972
rect 4567 1970 4576 1972
rect 4567 1961 4726 1970
rect 4567 1960 4576 1961
rect 4405 1913 4414 1940
rect 4536 1928 4545 1951
rect 4599 1952 4607 1961
rect 4676 1950 4682 1961
rect 4619 1929 4628 1940
rect 4323 1911 4344 1912
rect 4162 1893 4165 1899
rect 4201 1897 4204 1903
rect 4220 1897 4223 1903
rect 4230 1903 4233 1909
rect 4247 1903 4250 1909
rect 4323 1905 4370 1911
rect 4378 1906 4379 1911
rect 4323 1903 4371 1905
rect 4470 1921 4524 1925
rect 4536 1923 4578 1928
rect 4619 1923 4659 1929
rect 4230 1900 4250 1903
rect 4342 1899 4371 1903
rect 4186 1894 4257 1897
rect 4186 1893 4189 1894
rect 4161 1890 4189 1893
rect 4425 1891 4434 1901
rect 4470 1891 4477 1921
rect 4536 1920 4545 1923
rect 4619 1920 4628 1923
rect 4410 1884 4413 1888
rect 4425 1886 4477 1891
rect 4425 1877 4434 1886
rect 4486 1881 4490 1885
rect 4516 1888 4525 1908
rect 4597 1888 4606 1908
rect 4654 1911 4659 1923
rect 4689 1914 4700 1938
rect 4654 1906 4680 1911
rect 4689 1906 4715 1914
rect 4609 1899 4611 1903
rect 4689 1894 4700 1906
rect 3974 1856 4139 1859
rect 4405 1858 4413 1871
rect 4496 1858 4504 1876
rect 4579 1858 4587 1876
rect 4675 1858 4682 1888
rect 3336 1825 3657 1835
rect 3334 1804 3400 1813
rect 3456 1806 3535 1807
rect 3344 1778 3352 1804
rect 3392 1796 3400 1804
rect 3448 1798 3535 1806
rect 3448 1796 3456 1798
rect 3392 1787 3456 1796
rect 3475 1789 3483 1798
rect 3526 1796 3535 1798
rect 3526 1787 3685 1796
rect 3526 1786 3535 1787
rect 3364 1739 3373 1766
rect 3495 1754 3504 1777
rect 3558 1778 3566 1787
rect 3635 1776 3641 1787
rect 3757 1777 3872 1779
rect 3757 1776 3926 1777
rect 3578 1755 3587 1766
rect 3429 1747 3483 1751
rect 3495 1749 3537 1754
rect 3578 1749 3618 1755
rect 3384 1717 3393 1727
rect 3429 1717 3436 1747
rect 3495 1746 3504 1749
rect 3578 1746 3587 1749
rect 3369 1710 3372 1714
rect 3384 1712 3436 1717
rect 3384 1703 3393 1712
rect 3445 1707 3449 1711
rect 3475 1714 3484 1734
rect 3556 1714 3565 1734
rect 3613 1737 3618 1749
rect 3648 1740 3659 1764
rect 3757 1742 3760 1776
rect 3869 1774 3926 1776
rect 3770 1768 3798 1771
rect 3771 1762 3774 1768
rect 3795 1767 3798 1768
rect 3795 1764 3853 1767
rect 3858 1764 3866 1767
rect 3736 1741 3750 1742
rect 3736 1740 3757 1741
rect 3648 1738 3757 1740
rect 3613 1732 3639 1737
rect 3648 1733 3749 1738
rect 3762 1739 3772 1742
rect 3780 1742 3783 1750
rect 3810 1758 3813 1764
rect 3829 1758 3832 1764
rect 3780 1739 3801 1742
rect 3780 1736 3783 1739
rect 3648 1732 3674 1733
rect 3568 1725 3570 1729
rect 3648 1720 3659 1732
rect 3771 1726 3774 1730
rect 3765 1724 3789 1726
rect 3765 1723 3783 1724
rect 3788 1723 3789 1724
rect 3798 1716 3801 1739
rect 3839 1758 3859 1761
rect 3839 1752 3842 1758
rect 3856 1752 3859 1758
rect 3820 1731 3823 1734
rect 3820 1728 3838 1731
rect 3848 1721 3851 1728
rect 3869 1727 3872 1774
rect 3879 1765 3893 1768
rect 3898 1765 3913 1768
rect 3885 1759 3888 1765
rect 3869 1724 3896 1727
rect 3904 1726 3907 1735
rect 3904 1723 3910 1726
rect 3848 1718 3865 1721
rect 3770 1715 3789 1716
rect 3364 1684 3372 1697
rect 3455 1684 3463 1702
rect 3538 1684 3546 1702
rect 3634 1684 3641 1714
rect 3765 1713 3789 1715
rect 3798 1713 3841 1716
rect 3771 1707 3774 1713
rect 3827 1702 3852 1705
rect 3827 1700 3830 1702
rect 3726 1687 3753 1688
rect 3726 1684 3757 1687
rect 3337 1674 3658 1684
rect 3340 1649 3406 1658
rect 3462 1651 3541 1652
rect 3350 1623 3358 1649
rect 3398 1641 3406 1649
rect 3454 1643 3541 1651
rect 3454 1641 3462 1643
rect 3398 1632 3462 1641
rect 3481 1634 3489 1643
rect 3532 1641 3541 1643
rect 3532 1632 3691 1641
rect 3532 1631 3541 1632
rect 3370 1584 3379 1611
rect 3501 1599 3510 1622
rect 3564 1623 3572 1632
rect 3641 1621 3647 1632
rect 3584 1600 3593 1611
rect 3435 1592 3489 1596
rect 3501 1594 3543 1599
rect 3584 1594 3624 1600
rect 3390 1562 3399 1572
rect 3435 1562 3442 1592
rect 3501 1591 3510 1594
rect 3584 1591 3593 1594
rect 3375 1555 3378 1559
rect 3390 1557 3442 1562
rect 3390 1548 3399 1557
rect 3451 1552 3455 1556
rect 3481 1559 3490 1579
rect 3562 1559 3571 1579
rect 3619 1582 3624 1594
rect 3654 1585 3665 1609
rect 3726 1585 3743 1684
rect 3762 1684 3772 1687
rect 3780 1687 3783 1695
rect 3792 1697 3830 1700
rect 3862 1699 3865 1718
rect 3873 1718 3886 1721
rect 3792 1687 3795 1697
rect 3833 1696 3865 1699
rect 3833 1693 3836 1696
rect 3780 1684 3795 1687
rect 3759 1665 3762 1683
rect 3780 1681 3783 1684
rect 3832 1690 3838 1693
rect 3771 1671 3774 1675
rect 3792 1674 3797 1677
rect 3810 1677 3813 1681
rect 3857 1679 3860 1681
rect 3857 1677 3858 1679
rect 3802 1674 3858 1677
rect 3863 1674 3866 1677
rect 3792 1671 3795 1674
rect 3765 1668 3795 1671
rect 3873 1670 3876 1718
rect 3904 1720 3907 1723
rect 3895 1717 3907 1720
rect 3895 1714 3898 1717
rect 3885 1702 3888 1708
rect 3904 1702 3907 1708
rect 3923 1707 3926 1774
rect 3974 1759 3977 1856
rect 4378 1848 4699 1858
rect 4016 1794 4020 1797
rect 4025 1794 4056 1797
rect 4022 1788 4025 1794
rect 3971 1756 3977 1759
rect 4010 1753 4033 1756
rect 4041 1755 4044 1764
rect 4053 1766 4056 1794
rect 4081 1793 4118 1796
rect 4087 1787 4090 1793
rect 4115 1785 4118 1793
rect 4120 1780 4139 1783
rect 4078 1769 4098 1772
rect 4106 1767 4109 1775
rect 4121 1776 4124 1780
rect 4130 1767 4133 1770
rect 4053 1763 4061 1766
rect 4041 1752 4048 1755
rect 4016 1747 4023 1750
rect 4016 1737 4019 1747
rect 4041 1749 4044 1752
rect 4032 1746 4044 1749
rect 4032 1743 4035 1746
rect 3929 1733 3963 1736
rect 4010 1734 4019 1737
rect 3935 1727 3938 1733
rect 3954 1727 3957 1733
rect 4010 1732 4013 1734
rect 3971 1729 3989 1732
rect 3994 1729 4013 1732
rect 4022 1731 4025 1737
rect 4041 1731 4044 1737
rect 4058 1734 4061 1763
rect 4074 1763 4088 1766
rect 4074 1753 4077 1763
rect 4106 1764 4122 1767
rect 4106 1761 4109 1764
rect 4130 1764 4142 1767
rect 4096 1758 4109 1761
rect 4096 1755 4099 1758
rect 4130 1756 4133 1764
rect 4069 1750 4077 1753
rect 4087 1737 4090 1743
rect 4106 1737 4109 1743
rect 4121 1738 4124 1744
rect 4143 1738 4187 1741
rect 4115 1737 4146 1738
rect 4081 1735 4146 1737
rect 4081 1734 4139 1735
rect 4058 1731 4129 1734
rect 4156 1732 4159 1738
rect 4010 1723 4013 1729
rect 4016 1726 4046 1731
rect 4010 1720 4019 1723
rect 3944 1712 3947 1715
rect 3944 1709 3957 1712
rect 3923 1704 3936 1707
rect 3954 1706 3957 1709
rect 4016 1710 4019 1720
rect 4022 1720 4025 1726
rect 4041 1720 4044 1726
rect 4067 1725 4070 1731
rect 4101 1725 4104 1731
rect 4120 1725 4123 1731
rect 4032 1711 4035 1714
rect 4016 1707 4023 1710
rect 4032 1708 4044 1711
rect 3954 1703 3974 1706
rect 3879 1699 3916 1702
rect 3895 1693 3898 1699
rect 3919 1698 3946 1701
rect 3919 1670 3922 1698
rect 3954 1695 3957 1703
rect 3971 1695 3974 1703
rect 4041 1705 4044 1708
rect 4003 1701 4033 1704
rect 4041 1702 4068 1705
rect 4076 1705 4079 1713
rect 4110 1710 4113 1713
rect 4110 1707 4123 1710
rect 4184 1728 4187 1738
rect 4184 1725 4203 1728
rect 4233 1726 4261 1729
rect 4076 1702 4102 1705
rect 4120 1704 4123 1707
rect 3971 1692 3978 1695
rect 3983 1692 4010 1695
rect 4041 1693 4044 1702
rect 4076 1699 4079 1702
rect 4120 1701 4130 1704
rect 3935 1679 3938 1683
rect 3929 1674 3931 1677
rect 3936 1677 3938 1679
rect 3936 1674 3963 1677
rect 3798 1667 3922 1670
rect 4095 1696 4112 1699
rect 4120 1693 4123 1701
rect 4067 1689 4070 1693
rect 4061 1686 4067 1689
rect 4072 1686 4095 1689
rect 4092 1675 4095 1686
rect 4127 1696 4130 1701
rect 4146 1697 4167 1700
rect 4175 1699 4178 1708
rect 4190 1719 4193 1725
rect 4234 1720 4237 1726
rect 4258 1725 4261 1726
rect 4385 1725 4451 1734
rect 4507 1727 4586 1728
rect 4258 1722 4329 1725
rect 4175 1696 4191 1699
rect 4199 1699 4202 1707
rect 4199 1696 4220 1699
rect 4132 1691 4157 1694
rect 4175 1693 4178 1696
rect 4199 1693 4202 1696
rect 4225 1697 4235 1700
rect 4243 1700 4246 1708
rect 4273 1716 4276 1722
rect 4292 1716 4295 1722
rect 4243 1697 4264 1700
rect 4243 1694 4246 1697
rect 4166 1690 4178 1693
rect 4166 1687 4169 1690
rect 4190 1683 4193 1687
rect 4234 1684 4237 1688
rect 4208 1683 4252 1684
rect 4101 1675 4104 1681
rect 4156 1675 4159 1681
rect 4175 1675 4178 1681
rect 4184 1682 4252 1683
rect 4184 1681 4246 1682
rect 4184 1680 4211 1681
rect 4184 1675 4187 1680
rect 4092 1672 4113 1675
rect 4118 1672 4187 1675
rect 4251 1681 4252 1682
rect 4261 1674 4264 1697
rect 4302 1716 4322 1719
rect 4302 1710 4305 1716
rect 4319 1710 4322 1716
rect 4283 1689 4286 1692
rect 4283 1686 4301 1689
rect 4395 1699 4403 1725
rect 4443 1717 4451 1725
rect 4499 1719 4586 1727
rect 4499 1717 4507 1719
rect 4443 1708 4507 1717
rect 4526 1710 4534 1719
rect 4577 1717 4586 1719
rect 4577 1708 4736 1717
rect 4577 1707 4586 1708
rect 4311 1679 4314 1686
rect 4311 1676 4328 1679
rect 4233 1673 4252 1674
rect 4228 1671 4252 1673
rect 4261 1671 4304 1674
rect 3798 1665 3801 1667
rect 3759 1662 3801 1665
rect 4022 1663 4025 1669
rect 4234 1665 4237 1671
rect 4325 1665 4328 1676
rect 4016 1660 4020 1663
rect 4025 1660 4050 1663
rect 4325 1664 4329 1665
rect 4333 1664 4367 1665
rect 4290 1660 4315 1663
rect 4325 1661 4367 1664
rect 4290 1658 4293 1660
rect 4196 1642 4220 1645
rect 4196 1628 4199 1642
rect 4225 1642 4235 1645
rect 4243 1645 4246 1653
rect 4255 1655 4293 1658
rect 4325 1657 4328 1661
rect 4255 1645 4258 1655
rect 4296 1654 4328 1657
rect 4363 1659 4367 1661
rect 4415 1660 4424 1687
rect 4546 1675 4555 1698
rect 4609 1699 4617 1708
rect 4686 1697 4692 1708
rect 4629 1676 4638 1687
rect 4363 1658 4383 1659
rect 4363 1654 4379 1658
rect 4296 1651 4299 1654
rect 4363 1653 4367 1654
rect 4480 1668 4534 1672
rect 4546 1670 4588 1675
rect 4629 1670 4669 1676
rect 4243 1642 4258 1645
rect 4243 1639 4246 1642
rect 4295 1648 4301 1651
rect 4234 1629 4237 1633
rect 4255 1632 4260 1635
rect 4273 1635 4276 1639
rect 4320 1635 4323 1639
rect 4435 1638 4444 1648
rect 4480 1638 4487 1668
rect 4546 1667 4555 1670
rect 4629 1667 4638 1670
rect 4265 1632 4329 1635
rect 4255 1629 4258 1632
rect 4420 1631 4423 1635
rect 4435 1633 4487 1638
rect 3974 1625 4199 1628
rect 4228 1626 4258 1629
rect 3619 1577 3645 1582
rect 3654 1577 3744 1585
rect 3574 1570 3576 1574
rect 3654 1565 3665 1577
rect 3680 1576 3744 1577
rect 3370 1529 3378 1542
rect 3461 1529 3469 1547
rect 3544 1529 3552 1547
rect 3640 1529 3647 1559
rect 3757 1558 3872 1560
rect 3757 1557 3926 1558
rect 3343 1519 3664 1529
rect 3757 1523 3760 1557
rect 3869 1555 3926 1557
rect 3770 1549 3798 1552
rect 3771 1543 3774 1549
rect 3795 1548 3798 1549
rect 3795 1545 3853 1548
rect 3858 1545 3866 1548
rect 3705 1519 3757 1522
rect 3330 1502 3396 1511
rect 3452 1504 3531 1505
rect 3340 1476 3348 1502
rect 3388 1494 3396 1502
rect 3444 1496 3531 1504
rect 3444 1494 3452 1496
rect 3388 1485 3452 1494
rect 3471 1487 3479 1496
rect 3522 1494 3531 1496
rect 3522 1485 3681 1494
rect 3522 1484 3531 1485
rect 3360 1437 3369 1464
rect 3491 1452 3500 1475
rect 3554 1476 3562 1485
rect 3631 1474 3637 1485
rect 3574 1453 3583 1464
rect 3425 1445 3479 1449
rect 3491 1447 3533 1452
rect 3574 1447 3614 1453
rect 3380 1415 3389 1425
rect 3425 1415 3432 1445
rect 3491 1444 3500 1447
rect 3574 1444 3583 1447
rect 3365 1408 3368 1412
rect 3380 1410 3432 1415
rect 3380 1401 3389 1410
rect 3441 1405 3445 1409
rect 3471 1412 3480 1432
rect 3552 1412 3561 1432
rect 3609 1435 3614 1447
rect 3644 1438 3655 1462
rect 3705 1438 3717 1519
rect 3762 1520 3772 1523
rect 3780 1523 3783 1531
rect 3810 1539 3813 1545
rect 3829 1539 3832 1545
rect 3780 1520 3801 1523
rect 3780 1517 3783 1520
rect 3771 1507 3774 1511
rect 3765 1505 3789 1507
rect 3765 1504 3783 1505
rect 3788 1504 3789 1505
rect 3798 1497 3801 1520
rect 3839 1539 3859 1542
rect 3839 1533 3842 1539
rect 3856 1533 3859 1539
rect 3820 1512 3823 1515
rect 3820 1509 3838 1512
rect 3848 1502 3851 1509
rect 3869 1508 3872 1555
rect 3879 1546 3893 1549
rect 3898 1546 3913 1549
rect 3885 1540 3888 1546
rect 3869 1505 3896 1508
rect 3904 1507 3907 1516
rect 3904 1504 3910 1507
rect 3848 1499 3865 1502
rect 3770 1496 3789 1497
rect 3765 1494 3789 1496
rect 3798 1494 3841 1497
rect 3771 1488 3774 1494
rect 3827 1483 3852 1486
rect 3827 1481 3830 1483
rect 3609 1430 3635 1435
rect 3644 1430 3717 1438
rect 3731 1465 3757 1468
rect 3564 1423 3566 1427
rect 3644 1418 3655 1430
rect 3360 1382 3368 1395
rect 3451 1382 3459 1400
rect 3534 1382 3542 1400
rect 3630 1382 3637 1412
rect 3731 1385 3742 1465
rect 3762 1465 3772 1468
rect 3780 1468 3783 1476
rect 3792 1478 3830 1481
rect 3862 1480 3865 1499
rect 3873 1499 3886 1502
rect 3792 1468 3795 1478
rect 3833 1477 3865 1480
rect 3833 1474 3836 1477
rect 3780 1465 3795 1468
rect 3759 1446 3762 1464
rect 3780 1462 3783 1465
rect 3832 1471 3838 1474
rect 3771 1452 3774 1456
rect 3792 1455 3797 1458
rect 3810 1458 3813 1462
rect 3857 1460 3860 1462
rect 3857 1458 3858 1460
rect 3802 1455 3858 1458
rect 3863 1455 3866 1458
rect 3792 1452 3795 1455
rect 3765 1449 3795 1452
rect 3873 1451 3876 1499
rect 3904 1501 3907 1504
rect 3895 1498 3907 1501
rect 3895 1495 3898 1498
rect 3885 1483 3888 1489
rect 3904 1483 3907 1489
rect 3923 1488 3926 1555
rect 3974 1540 3977 1625
rect 4435 1624 4444 1633
rect 4496 1628 4500 1632
rect 4526 1635 4535 1655
rect 4607 1635 4616 1655
rect 4664 1658 4669 1670
rect 4699 1661 4710 1685
rect 4664 1653 4690 1658
rect 4699 1653 4725 1661
rect 4619 1646 4621 1650
rect 4699 1641 4710 1653
rect 4415 1605 4423 1618
rect 4506 1605 4514 1623
rect 4589 1605 4597 1623
rect 4685 1605 4692 1635
rect 4388 1595 4709 1605
rect 4016 1575 4020 1578
rect 4025 1575 4056 1578
rect 4022 1569 4025 1575
rect 3971 1537 3977 1540
rect 3996 1534 4033 1537
rect 4041 1536 4044 1545
rect 4053 1547 4056 1575
rect 4077 1574 4114 1577
rect 4083 1568 4086 1574
rect 4111 1566 4114 1574
rect 4116 1561 4135 1564
rect 4070 1550 4094 1553
rect 4102 1548 4105 1556
rect 4117 1557 4120 1561
rect 4126 1548 4129 1551
rect 4053 1544 4061 1547
rect 4041 1533 4048 1536
rect 4016 1528 4023 1531
rect 4016 1518 4019 1528
rect 4041 1530 4044 1533
rect 4032 1527 4044 1530
rect 4032 1524 4035 1527
rect 3929 1514 3963 1517
rect 4010 1515 4019 1518
rect 3935 1508 3938 1514
rect 3954 1508 3957 1514
rect 4010 1513 4013 1515
rect 3971 1510 4001 1513
rect 4006 1510 4013 1513
rect 4022 1512 4025 1518
rect 4041 1512 4044 1518
rect 4058 1515 4061 1544
rect 4072 1544 4084 1547
rect 4072 1534 4075 1544
rect 4102 1545 4118 1548
rect 4102 1542 4105 1545
rect 4126 1545 4137 1548
rect 4092 1539 4105 1542
rect 4092 1536 4095 1539
rect 4126 1537 4129 1545
rect 4069 1531 4075 1534
rect 4083 1518 4086 1524
rect 4102 1518 4105 1524
rect 4117 1519 4120 1525
rect 4143 1519 4186 1522
rect 4111 1518 4146 1519
rect 4077 1516 4146 1518
rect 4077 1515 4135 1516
rect 4058 1512 4129 1515
rect 4155 1513 4158 1519
rect 4010 1504 4013 1510
rect 4016 1507 4046 1512
rect 4010 1501 4019 1504
rect 3944 1493 3947 1496
rect 3944 1490 3957 1493
rect 3923 1485 3936 1488
rect 3954 1487 3957 1490
rect 4016 1491 4019 1501
rect 4022 1501 4025 1507
rect 4041 1501 4044 1507
rect 4067 1506 4070 1512
rect 4101 1506 4104 1512
rect 4120 1506 4123 1512
rect 4032 1492 4035 1495
rect 4016 1488 4023 1491
rect 4032 1489 4044 1492
rect 3954 1484 3974 1487
rect 3879 1480 3916 1483
rect 3895 1474 3898 1480
rect 3919 1479 3946 1482
rect 3919 1451 3922 1479
rect 3954 1476 3957 1484
rect 3971 1476 3974 1484
rect 4041 1486 4044 1489
rect 3982 1482 4033 1485
rect 4041 1483 4068 1486
rect 4076 1486 4079 1494
rect 4110 1491 4113 1494
rect 4110 1488 4123 1491
rect 4183 1509 4186 1519
rect 4385 1512 4451 1521
rect 4507 1514 4586 1515
rect 4183 1506 4202 1509
rect 4230 1507 4258 1510
rect 4076 1483 4102 1486
rect 4120 1485 4123 1488
rect 3971 1473 3981 1476
rect 3986 1473 4010 1476
rect 4041 1474 4044 1483
rect 4076 1480 4079 1483
rect 4120 1482 4130 1485
rect 3935 1460 3938 1464
rect 3929 1455 3931 1458
rect 3936 1458 3938 1460
rect 3936 1455 3963 1458
rect 3798 1448 3922 1451
rect 4095 1477 4112 1480
rect 4120 1474 4123 1482
rect 4067 1470 4070 1474
rect 4061 1467 4067 1470
rect 4072 1467 4095 1470
rect 4092 1456 4095 1467
rect 4127 1475 4130 1482
rect 4143 1478 4166 1481
rect 4174 1480 4177 1489
rect 4189 1500 4192 1506
rect 4231 1501 4234 1507
rect 4255 1506 4258 1507
rect 4255 1503 4326 1506
rect 4174 1477 4190 1480
rect 4198 1480 4201 1488
rect 4198 1477 4217 1480
rect 4127 1472 4156 1475
rect 4174 1474 4177 1477
rect 4198 1474 4201 1477
rect 4222 1478 4232 1481
rect 4240 1481 4243 1489
rect 4270 1497 4273 1503
rect 4289 1497 4292 1503
rect 4240 1478 4261 1481
rect 4240 1475 4243 1478
rect 4165 1471 4177 1474
rect 4165 1468 4168 1471
rect 4189 1464 4192 1468
rect 4231 1465 4234 1469
rect 4207 1464 4249 1465
rect 4101 1456 4104 1462
rect 4092 1453 4111 1456
rect 4155 1456 4158 1462
rect 4174 1456 4177 1462
rect 4183 1463 4249 1464
rect 4183 1462 4243 1463
rect 4183 1461 4210 1462
rect 4183 1456 4186 1461
rect 4116 1453 4186 1456
rect 4248 1462 4249 1463
rect 4258 1455 4261 1478
rect 4299 1497 4319 1500
rect 4299 1491 4302 1497
rect 4316 1491 4319 1497
rect 4280 1470 4283 1473
rect 4280 1467 4298 1470
rect 4395 1486 4403 1512
rect 4443 1504 4451 1512
rect 4499 1506 4586 1514
rect 4499 1504 4507 1506
rect 4443 1495 4507 1504
rect 4526 1497 4534 1506
rect 4577 1504 4586 1506
rect 4577 1495 4736 1504
rect 4577 1494 4586 1495
rect 4308 1460 4311 1467
rect 4308 1457 4325 1460
rect 4230 1454 4249 1455
rect 4225 1452 4249 1454
rect 4258 1452 4301 1455
rect 3798 1446 3801 1448
rect 3759 1443 3801 1446
rect 4022 1444 4025 1450
rect 4231 1446 4234 1452
rect 4322 1446 4325 1457
rect 4415 1447 4424 1474
rect 4546 1462 4555 1485
rect 4609 1486 4617 1495
rect 4686 1484 4692 1495
rect 4629 1463 4638 1474
rect 4016 1441 4020 1444
rect 4025 1441 4050 1444
rect 4322 1445 4326 1446
rect 4287 1441 4312 1444
rect 4322 1442 4379 1445
rect 4287 1439 4290 1441
rect 4197 1423 4217 1426
rect 4197 1404 4200 1423
rect 4222 1423 4232 1426
rect 4240 1426 4243 1434
rect 4252 1436 4290 1439
rect 4322 1438 4325 1442
rect 4330 1440 4379 1442
rect 4480 1455 4534 1459
rect 4546 1457 4588 1462
rect 4629 1457 4669 1463
rect 4252 1426 4255 1436
rect 4293 1435 4325 1438
rect 4293 1432 4296 1435
rect 4240 1423 4255 1426
rect 4240 1420 4243 1423
rect 4292 1429 4298 1432
rect 4435 1425 4444 1435
rect 4480 1425 4487 1455
rect 4546 1454 4555 1457
rect 4629 1454 4638 1457
rect 4231 1410 4234 1414
rect 4252 1413 4257 1416
rect 4270 1416 4273 1420
rect 4317 1416 4320 1420
rect 4420 1418 4423 1422
rect 4435 1420 4487 1425
rect 4262 1413 4326 1416
rect 4252 1410 4255 1413
rect 4435 1411 4444 1420
rect 4496 1415 4500 1419
rect 4526 1422 4535 1442
rect 4607 1422 4616 1442
rect 4664 1445 4669 1457
rect 4699 1448 4710 1472
rect 4664 1440 4690 1445
rect 4699 1440 4725 1448
rect 4619 1433 4621 1437
rect 4699 1428 4710 1440
rect 4225 1407 4255 1410
rect 3333 1372 3654 1382
rect 3693 1377 3742 1385
rect 3974 1401 4200 1404
rect 3331 1355 3397 1364
rect 3453 1357 3532 1358
rect 3341 1329 3349 1355
rect 3389 1347 3397 1355
rect 3445 1349 3532 1357
rect 3445 1347 3453 1349
rect 3389 1338 3453 1347
rect 3472 1340 3480 1349
rect 3523 1347 3532 1349
rect 3523 1338 3682 1347
rect 3523 1337 3532 1338
rect 3361 1290 3370 1317
rect 3492 1305 3501 1328
rect 3555 1329 3563 1338
rect 3632 1327 3638 1338
rect 3575 1306 3584 1317
rect 3426 1298 3480 1302
rect 3492 1300 3534 1305
rect 3575 1300 3615 1306
rect 3381 1268 3390 1278
rect 3426 1268 3433 1298
rect 3492 1297 3501 1300
rect 3575 1297 3584 1300
rect 3366 1261 3369 1265
rect 3381 1263 3433 1268
rect 3381 1254 3390 1263
rect 3442 1258 3446 1262
rect 3472 1265 3481 1285
rect 3553 1265 3562 1285
rect 3610 1288 3615 1300
rect 3645 1291 3656 1315
rect 3693 1291 3714 1377
rect 3757 1335 3872 1337
rect 3757 1334 3926 1335
rect 3757 1300 3760 1334
rect 3869 1332 3926 1334
rect 3770 1326 3798 1329
rect 3771 1320 3774 1326
rect 3795 1325 3798 1326
rect 3795 1322 3853 1325
rect 3858 1322 3866 1325
rect 3610 1283 3636 1288
rect 3645 1283 3714 1291
rect 3724 1296 3757 1299
rect 3565 1276 3567 1280
rect 3645 1271 3656 1283
rect 3361 1235 3369 1248
rect 3452 1235 3460 1253
rect 3535 1235 3543 1253
rect 3631 1235 3638 1265
rect 3334 1225 3655 1235
rect 3340 1193 3406 1202
rect 3462 1195 3541 1196
rect 3350 1167 3358 1193
rect 3398 1185 3406 1193
rect 3454 1187 3541 1195
rect 3454 1185 3462 1187
rect 3398 1176 3462 1185
rect 3481 1178 3489 1187
rect 3532 1185 3541 1187
rect 3532 1176 3691 1185
rect 3532 1175 3541 1176
rect 3370 1128 3379 1155
rect 3501 1143 3510 1166
rect 3564 1167 3572 1176
rect 3641 1165 3647 1176
rect 3584 1144 3593 1155
rect 3435 1136 3489 1140
rect 3501 1138 3543 1143
rect 3584 1138 3624 1144
rect 3390 1106 3399 1116
rect 3435 1106 3442 1136
rect 3501 1135 3510 1138
rect 3584 1135 3593 1138
rect 3375 1099 3378 1103
rect 3390 1101 3442 1106
rect 3390 1092 3399 1101
rect 3451 1096 3455 1100
rect 3481 1103 3490 1123
rect 3562 1103 3571 1123
rect 3619 1126 3624 1138
rect 3654 1129 3665 1153
rect 3724 1129 3729 1296
rect 3762 1297 3772 1300
rect 3780 1300 3783 1308
rect 3810 1316 3813 1322
rect 3829 1316 3832 1322
rect 3780 1297 3801 1300
rect 3780 1294 3783 1297
rect 3771 1284 3774 1288
rect 3765 1282 3789 1284
rect 3765 1281 3783 1282
rect 3788 1281 3789 1282
rect 3798 1274 3801 1297
rect 3839 1316 3859 1319
rect 3839 1310 3842 1316
rect 3856 1310 3859 1316
rect 3820 1289 3823 1292
rect 3820 1286 3838 1289
rect 3848 1279 3851 1286
rect 3869 1285 3872 1332
rect 3879 1323 3893 1326
rect 3898 1323 3913 1326
rect 3885 1317 3888 1323
rect 3869 1282 3896 1285
rect 3904 1284 3907 1293
rect 3904 1281 3910 1284
rect 3848 1276 3865 1279
rect 3770 1273 3789 1274
rect 3765 1271 3789 1273
rect 3798 1271 3841 1274
rect 3771 1265 3774 1271
rect 3827 1260 3852 1263
rect 3827 1258 3830 1260
rect 3619 1121 3645 1126
rect 3654 1123 3729 1129
rect 3743 1242 3757 1245
rect 3654 1121 3680 1123
rect 3574 1114 3576 1118
rect 3654 1109 3665 1121
rect 3370 1073 3378 1086
rect 3461 1073 3469 1091
rect 3544 1073 3552 1091
rect 3640 1073 3647 1103
rect 3343 1065 3664 1073
rect 3443 1063 3664 1065
rect 3343 1055 3408 1062
rect 3464 1057 3543 1058
rect 3352 1029 3360 1055
rect 3400 1047 3408 1055
rect 3456 1049 3543 1057
rect 3456 1047 3464 1049
rect 3400 1038 3464 1047
rect 3483 1040 3491 1049
rect 3534 1047 3543 1049
rect 3534 1038 3693 1047
rect 3534 1037 3543 1038
rect 3372 990 3381 1017
rect 3503 1005 3512 1028
rect 3566 1029 3574 1038
rect 3643 1027 3649 1038
rect 3586 1006 3595 1017
rect 3437 998 3491 1002
rect 3503 1000 3545 1005
rect 3586 1000 3626 1006
rect 3392 968 3401 978
rect 3437 968 3444 998
rect 3503 997 3512 1000
rect 3586 997 3595 1000
rect 3377 961 3380 965
rect 3392 963 3444 968
rect 3392 954 3401 963
rect 3453 958 3457 962
rect 3483 965 3492 985
rect 3564 965 3573 985
rect 3621 988 3626 1000
rect 3656 991 3667 1015
rect 3743 991 3750 1242
rect 3762 1242 3772 1245
rect 3780 1245 3783 1253
rect 3792 1255 3830 1258
rect 3862 1257 3865 1276
rect 3873 1276 3886 1279
rect 3792 1245 3795 1255
rect 3833 1254 3865 1257
rect 3833 1251 3836 1254
rect 3780 1242 3795 1245
rect 3759 1223 3762 1241
rect 3780 1239 3783 1242
rect 3832 1248 3838 1251
rect 3771 1229 3774 1233
rect 3792 1232 3797 1235
rect 3810 1235 3813 1239
rect 3857 1237 3860 1239
rect 3857 1235 3858 1237
rect 3802 1232 3858 1235
rect 3863 1232 3866 1235
rect 3792 1229 3795 1232
rect 3765 1226 3795 1229
rect 3873 1228 3876 1276
rect 3904 1278 3907 1281
rect 3895 1275 3907 1278
rect 3895 1272 3898 1275
rect 3885 1260 3888 1266
rect 3904 1260 3907 1266
rect 3923 1265 3926 1332
rect 3974 1317 3977 1401
rect 4415 1392 4423 1405
rect 4506 1392 4514 1410
rect 4589 1392 4597 1410
rect 4685 1392 4692 1422
rect 4388 1382 4709 1392
rect 4013 1352 4017 1355
rect 4133 1355 4190 1358
rect 4022 1352 4053 1355
rect 4019 1346 4022 1352
rect 3971 1314 3977 1317
rect 4006 1311 4030 1314
rect 4038 1313 4041 1322
rect 4050 1324 4053 1352
rect 4075 1351 4112 1354
rect 4081 1345 4084 1351
rect 4109 1343 4112 1351
rect 4133 1341 4136 1355
rect 4114 1338 4136 1341
rect 4159 1349 4162 1355
rect 4070 1327 4092 1330
rect 4100 1325 4103 1333
rect 4115 1334 4118 1338
rect 4187 1345 4190 1355
rect 4217 1356 4257 1359
rect 4217 1345 4220 1356
rect 4187 1342 4220 1345
rect 4226 1350 4229 1356
rect 4150 1331 4170 1334
rect 4178 1329 4181 1337
rect 4193 1338 4196 1342
rect 4254 1346 4257 1356
rect 4254 1343 4278 1346
rect 4220 1332 4237 1335
rect 4202 1329 4205 1332
rect 4245 1330 4248 1338
rect 4260 1339 4263 1343
rect 4269 1330 4272 1333
rect 4124 1325 4127 1328
rect 4147 1327 4160 1328
rect 4050 1321 4058 1324
rect 4038 1310 4045 1313
rect 4013 1305 4020 1308
rect 4013 1295 4016 1305
rect 4038 1307 4041 1310
rect 4029 1304 4041 1307
rect 4029 1301 4032 1304
rect 3929 1291 3963 1294
rect 4007 1292 4016 1295
rect 3935 1285 3938 1291
rect 3954 1285 3957 1291
rect 4007 1290 4010 1292
rect 3971 1287 4010 1290
rect 4019 1289 4022 1295
rect 4038 1289 4041 1295
rect 4055 1292 4058 1321
rect 4069 1321 4082 1324
rect 4069 1311 4072 1321
rect 4100 1322 4116 1325
rect 4100 1319 4103 1322
rect 4124 1322 4131 1325
rect 4150 1325 4160 1327
rect 4178 1326 4194 1329
rect 4178 1323 4181 1326
rect 4202 1326 4227 1329
rect 4090 1316 4103 1319
rect 4090 1313 4093 1316
rect 4124 1314 4127 1322
rect 4168 1320 4181 1323
rect 4168 1317 4171 1320
rect 4202 1318 4205 1326
rect 4245 1327 4261 1330
rect 4245 1324 4248 1327
rect 4269 1327 4275 1330
rect 4235 1321 4248 1324
rect 4235 1318 4238 1321
rect 4269 1319 4272 1327
rect 4382 1322 4448 1331
rect 4504 1324 4583 1325
rect 4066 1308 4072 1311
rect 4081 1295 4084 1301
rect 4100 1295 4103 1301
rect 4115 1296 4118 1302
rect 4159 1299 4162 1305
rect 4178 1299 4181 1305
rect 4193 1300 4196 1306
rect 4226 1300 4229 1306
rect 4245 1300 4248 1306
rect 4260 1301 4263 1307
rect 4254 1300 4278 1301
rect 4187 1299 4278 1300
rect 4153 1298 4278 1299
rect 4153 1297 4257 1298
rect 4153 1296 4190 1297
rect 4392 1296 4400 1322
rect 4440 1314 4448 1322
rect 4496 1316 4583 1324
rect 4496 1314 4504 1316
rect 4440 1305 4504 1314
rect 4523 1307 4531 1316
rect 4574 1314 4583 1316
rect 4574 1305 4733 1314
rect 4574 1304 4583 1305
rect 4109 1295 4177 1296
rect 4075 1293 4177 1295
rect 4075 1292 4133 1293
rect 4055 1289 4126 1292
rect 4007 1281 4010 1287
rect 4013 1284 4043 1289
rect 4007 1278 4016 1281
rect 3944 1270 3947 1273
rect 3944 1267 3957 1270
rect 3923 1262 3936 1265
rect 3954 1264 3957 1267
rect 4013 1268 4016 1278
rect 4019 1278 4022 1284
rect 4038 1278 4041 1284
rect 4064 1283 4067 1289
rect 4098 1283 4101 1289
rect 4117 1283 4120 1289
rect 4029 1269 4032 1272
rect 4146 1287 4149 1293
rect 4013 1265 4020 1268
rect 4029 1266 4041 1269
rect 3954 1261 3974 1264
rect 3879 1257 3916 1260
rect 3895 1251 3898 1257
rect 3919 1256 3946 1259
rect 3919 1228 3922 1256
rect 3954 1253 3957 1261
rect 3971 1253 3974 1261
rect 4038 1263 4041 1266
rect 3986 1259 4030 1262
rect 4038 1260 4065 1263
rect 4073 1263 4076 1271
rect 4107 1268 4110 1271
rect 4107 1265 4120 1268
rect 4073 1260 4099 1263
rect 4117 1262 4120 1265
rect 4174 1283 4177 1293
rect 4174 1280 4244 1283
rect 3971 1250 4007 1253
rect 4038 1251 4041 1260
rect 4073 1257 4076 1260
rect 4117 1259 4127 1262
rect 3935 1237 3938 1241
rect 3929 1232 3931 1235
rect 3936 1235 3938 1237
rect 3936 1232 3963 1235
rect 3798 1225 3922 1228
rect 4092 1254 4109 1257
rect 4117 1251 4120 1259
rect 4064 1247 4067 1251
rect 4058 1244 4064 1247
rect 4069 1244 4092 1247
rect 4089 1233 4092 1244
rect 4124 1249 4127 1259
rect 4136 1252 4157 1255
rect 4165 1254 4168 1263
rect 4180 1274 4183 1280
rect 4213 1274 4216 1280
rect 4165 1251 4181 1254
rect 4189 1254 4192 1262
rect 4189 1251 4204 1254
rect 4124 1246 4147 1249
rect 4165 1248 4168 1251
rect 4189 1248 4192 1251
rect 4156 1245 4168 1248
rect 4156 1242 4159 1245
rect 4201 1242 4204 1251
rect 4241 1270 4244 1280
rect 4241 1267 4265 1270
rect 4098 1233 4101 1239
rect 4180 1238 4183 1242
rect 4201 1239 4224 1242
rect 4232 1241 4235 1250
rect 4247 1261 4250 1267
rect 4232 1238 4248 1241
rect 4256 1241 4259 1249
rect 4284 1259 4371 1260
rect 4284 1256 4368 1259
rect 4284 1241 4287 1256
rect 4366 1252 4368 1256
rect 4412 1257 4421 1284
rect 4543 1272 4552 1295
rect 4606 1296 4614 1305
rect 4683 1294 4689 1305
rect 4626 1273 4635 1284
rect 4366 1251 4381 1252
rect 4477 1265 4531 1269
rect 4543 1267 4585 1272
rect 4626 1267 4666 1273
rect 4256 1238 4287 1241
rect 4089 1230 4107 1233
rect 4112 1230 4126 1233
rect 4146 1230 4149 1236
rect 4165 1230 4168 1236
rect 4174 1235 4198 1238
rect 4174 1230 4177 1235
rect 3798 1223 3801 1225
rect 3759 1220 3801 1223
rect 4019 1221 4022 1227
rect 4013 1218 4017 1221
rect 4022 1218 4047 1221
rect 4109 1207 4112 1230
rect 4123 1227 4177 1230
rect 4195 1217 4198 1235
rect 4207 1233 4214 1236
rect 4232 1235 4235 1238
rect 4256 1235 4259 1238
rect 4223 1232 4235 1235
rect 4223 1229 4226 1232
rect 4432 1235 4441 1245
rect 4477 1235 4484 1265
rect 4543 1264 4552 1267
rect 4626 1264 4635 1267
rect 4247 1225 4250 1229
rect 4417 1228 4420 1232
rect 4432 1230 4484 1235
rect 4213 1217 4216 1223
rect 4232 1217 4235 1223
rect 4241 1222 4265 1225
rect 4241 1217 4244 1222
rect 4432 1221 4441 1230
rect 4493 1225 4497 1229
rect 4523 1232 4532 1252
rect 4604 1232 4613 1252
rect 4661 1255 4666 1267
rect 4696 1258 4707 1282
rect 4661 1250 4687 1255
rect 4696 1250 4722 1258
rect 4616 1243 4618 1247
rect 4696 1238 4707 1250
rect 4195 1214 4244 1217
rect 3770 1204 3799 1207
rect 3804 1204 4301 1207
rect 4412 1202 4420 1215
rect 4503 1202 4511 1220
rect 4586 1202 4594 1220
rect 4682 1202 4689 1232
rect 4385 1192 4706 1202
rect 3621 983 3647 988
rect 3656 983 3750 991
rect 3576 976 3578 980
rect 3656 971 3667 983
rect 3682 982 3750 983
rect 3372 935 3380 948
rect 3463 935 3471 953
rect 3546 935 3554 953
rect 3642 935 3649 965
rect 3345 925 3666 935
<< m2contact >>
rect 4121 2147 4126 2152
rect 3974 2093 3979 2098
rect 3757 1978 3762 1983
rect 3757 1924 3762 1929
rect 3865 1944 3870 1949
rect 3910 1962 3915 1967
rect 4059 2108 4064 2113
rect 4028 2094 4033 2099
rect 4121 2093 4126 2098
rect 3966 1995 3971 2000
rect 4149 1989 4154 1994
rect 3966 1968 3971 1973
rect 4003 1968 4008 1973
rect 4077 1967 4082 1972
rect 4114 1973 4119 1978
rect 4148 1973 4153 1978
rect 3996 1943 4001 1948
rect 4067 1944 4072 1949
rect 4122 1945 4127 1950
rect 4148 1919 4153 1924
rect 3757 1737 3762 1742
rect 3757 1683 3762 1688
rect 3865 1703 3870 1708
rect 3910 1721 3915 1726
rect 4020 1794 4025 1799
rect 3966 1754 3971 1759
rect 4005 1753 4010 1758
rect 4073 1769 4078 1774
rect 3966 1727 3971 1732
rect 3989 1727 3994 1732
rect 4064 1750 4069 1755
rect 4142 1764 4147 1769
rect 4046 1726 4051 1731
rect 3998 1701 4003 1706
rect 3978 1691 3983 1696
rect 4067 1684 4072 1689
rect 4141 1697 4146 1702
rect 4127 1691 4132 1696
rect 4220 1695 4225 1700
rect 4020 1658 4025 1663
rect 4220 1641 4225 1646
rect 3757 1518 3762 1523
rect 3757 1464 3762 1469
rect 3865 1484 3870 1489
rect 3910 1502 3915 1507
rect 4020 1575 4025 1580
rect 3966 1535 3971 1540
rect 3991 1534 3996 1539
rect 4065 1550 4070 1555
rect 4048 1531 4053 1536
rect 3966 1508 3971 1513
rect 4001 1508 4006 1513
rect 4064 1531 4069 1536
rect 4137 1543 4142 1548
rect 4046 1507 4051 1512
rect 3977 1482 3982 1487
rect 3981 1471 3986 1476
rect 4067 1465 4072 1470
rect 4138 1478 4143 1483
rect 4217 1476 4222 1481
rect 4020 1439 4025 1444
rect 4217 1422 4222 1427
rect 3757 1295 3762 1300
rect 3757 1241 3762 1246
rect 3865 1261 3870 1266
rect 3910 1279 3915 1284
rect 4017 1352 4022 1357
rect 3966 1312 3971 1317
rect 4001 1311 4006 1316
rect 4109 1338 4114 1343
rect 4065 1327 4070 1332
rect 4045 1308 4050 1313
rect 3966 1285 3971 1290
rect 4131 1322 4136 1327
rect 4043 1284 4048 1289
rect 3981 1259 3986 1264
rect 4064 1242 4069 1247
rect 4131 1252 4136 1257
rect 4107 1230 4112 1235
rect 4017 1216 4022 1221
<< pm12contact >>
rect 3813 1961 3818 1966
rect 3822 1960 3827 1965
rect 4177 2110 4182 2115
rect 4186 2111 4191 2116
rect 4204 1936 4209 1941
rect 4213 1937 4218 1942
rect 3813 1720 3818 1725
rect 3822 1719 3827 1724
rect 4276 1678 4281 1683
rect 4285 1677 4290 1682
rect 3813 1501 3818 1506
rect 3822 1500 3827 1505
rect 4273 1459 4278 1464
rect 4282 1458 4287 1463
rect 3813 1278 3818 1283
rect 3822 1277 3827 1282
<< metal2 >>
rect 4123 2129 4126 2147
rect 4123 2126 4189 2129
rect 4186 2116 4189 2126
rect 4156 2110 4177 2113
rect 3979 2095 4028 2098
rect 3867 1997 3966 2000
rect 3758 1972 3761 1978
rect 3758 1969 3795 1972
rect 3792 1966 3795 1969
rect 3792 1963 3813 1966
rect 3822 1950 3825 1960
rect 3759 1947 3825 1950
rect 3867 1949 3870 1997
rect 3919 1970 3966 1973
rect 3919 1967 3922 1970
rect 3915 1964 3922 1967
rect 3759 1929 3762 1947
rect 3867 1756 3966 1759
rect 3758 1731 3761 1737
rect 3758 1728 3795 1731
rect 3792 1725 3795 1728
rect 3792 1722 3813 1725
rect 3822 1709 3825 1719
rect 3759 1706 3825 1709
rect 3867 1708 3870 1756
rect 3919 1729 3966 1732
rect 3919 1726 3922 1729
rect 3915 1723 3922 1726
rect 3759 1688 3762 1706
rect 3867 1537 3966 1540
rect 3758 1512 3761 1518
rect 3758 1509 3795 1512
rect 3792 1506 3795 1509
rect 3792 1503 3813 1506
rect 3822 1490 3825 1500
rect 3759 1487 3825 1490
rect 3867 1489 3870 1537
rect 3919 1510 3966 1513
rect 3919 1507 3922 1510
rect 3915 1504 3922 1507
rect 3759 1469 3762 1487
rect 3979 1487 3982 1691
rect 3991 1539 3994 1727
rect 3998 1706 4001 1943
rect 4005 1758 4008 1968
rect 4021 1799 4024 2020
rect 4020 1663 4023 1794
rect 4060 1772 4063 2108
rect 4156 2107 4159 2110
rect 4122 2104 4159 2107
rect 4122 2098 4125 2104
rect 4150 1994 4153 2052
rect 4124 1990 4149 1993
rect 4077 1949 4080 1967
rect 4072 1946 4080 1949
rect 4114 1805 4117 1973
rect 4124 1950 4127 1990
rect 4150 1955 4153 1973
rect 4150 1952 4216 1955
rect 4213 1942 4216 1952
rect 4183 1936 4204 1939
rect 4183 1933 4186 1936
rect 4149 1930 4186 1933
rect 4149 1924 4152 1930
rect 4103 1802 4117 1805
rect 4060 1769 4073 1772
rect 4053 1750 4064 1753
rect 4051 1726 4056 1729
rect 4053 1687 4056 1726
rect 4053 1684 4067 1687
rect 4021 1580 4024 1658
rect 4103 1635 4106 1802
rect 4142 1702 4145 1764
rect 4065 1632 4106 1635
rect 3867 1314 3966 1317
rect 3758 1289 3761 1295
rect 3758 1286 3795 1289
rect 3792 1283 3795 1286
rect 3792 1280 3813 1283
rect 3822 1267 3825 1277
rect 3759 1264 3825 1267
rect 3867 1266 3870 1314
rect 3919 1287 3966 1290
rect 3919 1284 3922 1287
rect 3915 1281 3922 1284
rect 3759 1246 3762 1264
rect 3983 1264 3986 1471
rect 4003 1316 4006 1508
rect 4020 1444 4023 1575
rect 4065 1555 4068 1632
rect 4129 1609 4132 1691
rect 4221 1689 4224 1695
rect 4221 1686 4258 1689
rect 4255 1683 4258 1686
rect 4255 1680 4276 1683
rect 4285 1667 4288 1677
rect 4222 1664 4288 1667
rect 4222 1646 4225 1664
rect 4081 1606 4132 1609
rect 4053 1531 4064 1534
rect 4051 1507 4056 1510
rect 4053 1468 4056 1507
rect 4053 1465 4067 1468
rect 4022 1435 4025 1439
rect 4019 1432 4025 1435
rect 4019 1357 4022 1432
rect 4081 1368 4084 1606
rect 4138 1483 4141 1543
rect 4218 1470 4221 1476
rect 4218 1467 4255 1470
rect 4252 1464 4255 1467
rect 4065 1365 4084 1368
rect 4252 1461 4273 1464
rect 4017 1221 4020 1352
rect 4065 1332 4068 1365
rect 4111 1343 4114 1453
rect 4282 1448 4285 1458
rect 4219 1445 4285 1448
rect 4219 1427 4222 1445
rect 4050 1308 4061 1311
rect 4048 1284 4053 1287
rect 4050 1245 4053 1284
rect 4050 1242 4064 1245
rect 4109 1235 4112 1338
rect 4131 1257 4134 1322
<< m123contact >>
rect 3893 2199 3898 2204
rect 4025 2199 4030 2204
rect 4129 2199 4134 2204
rect 4161 2156 4166 2161
rect 4101 2119 4106 2124
rect 4129 2115 4134 2120
rect 4147 2111 4152 2116
rect 3765 2009 3770 2014
rect 3853 2005 3858 2010
rect 3893 2006 3898 2011
rect 3765 1956 3770 1961
rect 3783 1960 3788 1965
rect 3938 1977 3943 1982
rect 3894 1929 3899 1934
rect 3797 1915 3802 1920
rect 3858 1915 3863 1920
rect 3931 1915 3936 1920
rect 3765 1768 3770 1773
rect 3853 1764 3858 1769
rect 3893 1765 3898 1770
rect 3765 1715 3770 1720
rect 3783 1719 3788 1724
rect 3938 1736 3943 1741
rect 3894 1688 3899 1693
rect 3797 1674 3802 1679
rect 3858 1674 3863 1679
rect 3931 1674 3936 1679
rect 3765 1549 3770 1554
rect 3853 1545 3858 1550
rect 3893 1546 3898 1551
rect 3765 1496 3770 1501
rect 3783 1500 3788 1505
rect 3938 1517 3943 1522
rect 4024 2017 4029 2022
rect 4010 1692 4015 1697
rect 4129 2062 4134 2067
rect 4149 2052 4154 2057
rect 4119 2003 4124 2008
rect 4101 1943 4106 1948
rect 4188 1982 4193 1987
rect 4156 1941 4161 1946
rect 4174 1937 4179 1942
rect 4156 1888 4161 1893
rect 4048 1750 4053 1755
rect 4090 1694 4095 1699
rect 4115 1780 4120 1785
rect 4203 1725 4208 1730
rect 4228 1726 4233 1731
rect 4113 1670 4118 1675
rect 3894 1469 3899 1474
rect 3797 1455 3802 1460
rect 3858 1455 3863 1460
rect 3931 1455 3936 1460
rect 3765 1326 3770 1331
rect 3853 1322 3858 1327
rect 3893 1323 3898 1328
rect 3765 1273 3770 1278
rect 3783 1277 3788 1282
rect 3938 1294 3943 1299
rect 4010 1473 4015 1478
rect 4228 1673 4233 1678
rect 4246 1677 4251 1682
rect 4260 1632 4265 1637
rect 4111 1561 4116 1566
rect 4202 1506 4207 1511
rect 4225 1507 4230 1512
rect 4090 1475 4095 1480
rect 4111 1453 4116 1458
rect 4225 1454 4230 1459
rect 4243 1458 4248 1463
rect 3894 1246 3899 1251
rect 4007 1250 4012 1255
rect 3797 1232 3802 1237
rect 3858 1232 3863 1237
rect 3931 1232 3936 1237
rect 4257 1413 4262 1418
rect 4061 1308 4066 1313
rect 4087 1252 4092 1257
rect 4145 1331 4150 1336
rect 4215 1332 4220 1337
rect 4275 1327 4280 1332
rect 4145 1322 4150 1327
rect 4202 1231 4207 1236
rect 3799 1202 3804 1207
<< metal3 >>
rect 3894 2011 3897 2199
rect 4026 2022 4029 2199
rect 4130 2120 4133 2199
rect 4103 2045 4106 2119
rect 4161 2116 4164 2156
rect 4129 2067 4132 2115
rect 4152 2113 4164 2116
rect 4149 2057 4152 2111
rect 4103 2042 4239 2045
rect 3765 1961 3768 2009
rect 3858 2007 3893 2010
rect 3898 2006 3919 2009
rect 3916 1980 3919 2006
rect 4124 2004 4136 2007
rect 3916 1977 3938 1980
rect 3788 1960 3800 1963
rect 3797 1920 3800 1960
rect 3802 1915 3809 1918
rect 3895 1918 3898 1929
rect 3863 1915 3931 1918
rect 3765 1720 3768 1768
rect 3788 1719 3800 1722
rect 3797 1679 3800 1719
rect 3806 1677 3809 1915
rect 3858 1766 3893 1769
rect 3898 1765 3919 1768
rect 3916 1739 3919 1765
rect 3916 1736 3938 1739
rect 3802 1674 3809 1677
rect 3895 1677 3898 1688
rect 3863 1674 3931 1677
rect 3765 1501 3768 1549
rect 3788 1500 3800 1503
rect 3797 1460 3800 1500
rect 3785 1456 3797 1459
rect 3765 1278 3768 1326
rect 3785 1282 3788 1456
rect 3806 1458 3809 1674
rect 3858 1547 3893 1550
rect 3898 1546 3919 1549
rect 3916 1520 3919 1546
rect 3916 1517 3938 1520
rect 3802 1455 3809 1458
rect 3895 1458 3898 1469
rect 3863 1455 3931 1458
rect 3858 1324 3893 1327
rect 3898 1323 3919 1326
rect 3916 1297 3919 1323
rect 3916 1294 3938 1297
rect 3943 1294 3946 1982
rect 4133 1946 4136 2004
rect 4133 1943 4156 1946
rect 4102 1824 4105 1943
rect 4188 1942 4191 1982
rect 4156 1893 4159 1941
rect 4179 1939 4191 1942
rect 4102 1821 4118 1824
rect 4115 1785 4118 1821
rect 4236 1789 4239 2042
rect 4236 1786 4311 1789
rect 4050 1707 4053 1750
rect 4050 1704 4102 1707
rect 4015 1694 4090 1697
rect 4015 1475 4090 1478
rect 4099 1374 4102 1704
rect 4115 1675 4118 1780
rect 4208 1727 4228 1730
rect 4228 1678 4231 1726
rect 4251 1677 4263 1680
rect 4113 1566 4116 1670
rect 4260 1637 4263 1677
rect 4112 1458 4115 1561
rect 4207 1507 4225 1510
rect 4225 1459 4228 1507
rect 4248 1458 4260 1461
rect 4257 1418 4260 1458
rect 4308 1385 4311 1786
rect 4215 1382 4311 1385
rect 4099 1371 4148 1374
rect 4145 1336 4148 1371
rect 4215 1337 4218 1382
rect 4145 1311 4148 1322
rect 4066 1308 4148 1311
rect 4280 1291 4283 1330
rect 4204 1288 4283 1291
rect 3788 1277 3800 1280
rect 3797 1237 3800 1277
rect 4012 1252 4087 1255
rect 3895 1235 3898 1246
rect 3863 1232 3931 1235
rect 4204 1236 4207 1288
rect 3799 1207 3802 1232
<< labels >>
rlabel metal1 4718 1253 4718 1253 1 cout
rlabel polysilicon 4383 1252 4383 1252 1 p5
rlabel metal1 4721 1443 4721 1443 1 s4
rlabel polycontact 4386 1442 4386 1442 1 p4
rlabel metal1 4721 1656 4721 1656 1 s3
rlabel polysilicon 4386 1655 4386 1655 1 p3
rlabel polycontact 4376 1908 4376 1908 1 p2
rlabel metal1 4711 1909 4711 1909 1 s2
rlabel metal1 4675 2108 4675 2108 1 s1
rlabel polysilicon 4340 2107 4340 2107 1 p1
rlabel polysilicon 3343 985 3343 985 1 y4
rlabel metal1 3678 986 3678 986 1 b4
rlabel polysilicon 3341 1123 3341 1123 1 x4
rlabel metal1 3676 1124 3676 1124 1 a4
rlabel metal1 3667 1286 3667 1286 1 b3
rlabel polysilicon 3332 1285 3332 1285 1 y3
rlabel metal1 3665 1433 3666 1433 1 a3
rlabel polysilicon 3331 1432 3331 1432 1 x3
rlabel metal1 3676 1580 3676 1580 1 b2
rlabel polysilicon 3341 1579 3341 1579 1 y2
rlabel metal1 3670 1735 3670 1735 1 a2
rlabel polysilicon 3335 1734 3335 1734 1 x2
rlabel metal1 3668 1886 3669 1886 1 b1
rlabel polysilicon 3334 1885 3334 1885 1 y1
rlabel metal1 3662 2039 3662 2039 1 a1
rlabel polysilicon 3327 2038 3327 2038 1 x1
rlabel metal1 4617 1244 4617 1244 1 clk
rlabel metal1 4496 1226 4496 1226 1 clk
rlabel metal1 4418 1230 4418 1230 1 clk
rlabel metal1 4526 1320 4526 1320 5 vdd
rlabel metal1 4506 1198 4506 1198 1 gnd
rlabel metal1 4620 1434 4620 1434 1 clk
rlabel metal1 4499 1416 4499 1416 1 clk
rlabel metal1 4421 1420 4421 1420 1 clk
rlabel metal1 4529 1510 4529 1510 5 vdd
rlabel metal1 4509 1388 4509 1388 1 gnd
rlabel metal1 4620 1647 4620 1647 1 clk
rlabel metal1 4499 1629 4499 1629 1 clk
rlabel metal1 4421 1633 4421 1633 1 clk
rlabel metal1 4529 1723 4529 1723 5 vdd
rlabel metal1 4509 1601 4509 1601 1 gnd
rlabel metal1 4610 1900 4610 1900 1 clk
rlabel metal1 4489 1882 4489 1882 1 clk
rlabel metal1 4411 1886 4411 1886 1 clk
rlabel metal1 4519 1976 4519 1976 5 vdd
rlabel metal1 4499 1854 4499 1854 1 gnd
rlabel metal1 4574 2099 4574 2099 1 clk
rlabel metal1 4453 2081 4453 2081 1 clk
rlabel metal1 4375 2085 4375 2085 1 clk
rlabel metal1 4483 2175 4483 2175 5 vdd
rlabel metal1 4463 2053 4463 2053 1 gnd
rlabel metal1 3577 977 3577 977 1 clk
rlabel metal1 3456 959 3456 959 1 clk
rlabel metal1 3378 963 3378 963 1 clk
rlabel metal1 3486 1053 3486 1053 5 vdd
rlabel metal1 3466 931 3466 931 1 gnd
rlabel metal1 3575 1115 3575 1115 1 clk
rlabel metal1 3454 1097 3454 1097 1 clk
rlabel metal1 3376 1101 3376 1101 1 clk
rlabel metal1 3484 1191 3484 1191 5 vdd
rlabel metal1 3464 1069 3464 1069 1 gnd
rlabel metal1 3566 1277 3566 1277 1 clk
rlabel metal1 3445 1259 3445 1259 1 clk
rlabel metal1 3367 1263 3367 1263 1 clk
rlabel metal1 3475 1353 3475 1353 5 vdd
rlabel metal1 3455 1231 3455 1231 1 gnd
rlabel metal1 3454 1378 3454 1378 1 gnd
rlabel metal1 3474 1500 3474 1500 5 vdd
rlabel metal1 3366 1410 3366 1410 1 clk
rlabel metal1 3444 1406 3444 1406 1 clk
rlabel metal1 3565 1424 3565 1424 1 clk
rlabel metal1 3575 1571 3575 1571 1 clk
rlabel metal1 3454 1553 3454 1553 1 clk
rlabel metal1 3376 1557 3376 1557 1 clk
rlabel metal1 3484 1647 3484 1647 5 vdd
rlabel metal1 3464 1525 3464 1525 1 gnd
rlabel metal1 3458 1680 3458 1680 1 gnd
rlabel metal1 3478 1802 3478 1802 5 vdd
rlabel metal1 3370 1712 3370 1712 1 clk
rlabel metal1 3448 1708 3448 1708 1 clk
rlabel metal1 3569 1726 3569 1726 1 clk
rlabel metal1 3568 1877 3568 1877 1 clk
rlabel metal1 3447 1859 3447 1859 1 clk
rlabel metal1 3369 1863 3369 1863 1 clk
rlabel metal1 3477 1953 3477 1953 5 vdd
rlabel metal1 3457 1831 3457 1831 1 gnd
rlabel metal1 3561 2030 3561 2030 1 clk
rlabel metal1 3440 2012 3440 2012 1 clk
rlabel metal1 3362 2016 3362 2016 1 clk
rlabel metal1 3470 2106 3470 2106 5 vdd
rlabel metal1 3450 1984 3450 1984 1 gnd
rlabel metal1 4149 2166 4149 2166 5 gnd!
rlabel metal1 4160 2160 4160 2160 5 gnd!
rlabel metal1 4199 2160 4199 2160 5 gnd!
rlabel metal1 4228 1216 4228 1216 1 gnd!
rlabel metal1 4031 1220 4031 1220 1 vdd!
rlabel metal1 3826 2175 3826 2178 1 cin
rlabel metal1 3813 1205 3813 1205 1 gnd!
rlabel metal1 3967 1206 3967 1206 1 gnd
rlabel metal1 3988 2200 3988 2200 5 vdd
<< end >>
