magic
tech scmos
timestamp 1731956492
<< metal1 >>
rect 29 90 38 93
rect 35 62 38 90
rect 35 59 43 62
rect -9 49 -2 52
rect -2 33 1 46
rect -8 30 1 33
rect -8 28 -5 30
rect -9 25 -5 28
rect 40 27 43 59
rect 51 46 52 49
rect 67 27 77 30
rect -8 19 -5 25
rect -8 16 1 19
rect -2 3 1 16
rect -9 -3 -2 0
rect 32 -2 43 1
rect 67 -2 77 1
rect 111 -3 112 0
rect -9 -12 -8 -9
rect 67 -18 77 -15
rect 74 -29 77 -18
rect 74 -32 82 -29
<< m2contact >>
rect 2 90 7 95
rect 30 46 35 51
rect 46 46 51 51
rect 28 22 33 27
rect 49 -20 54 -15
rect 2 -46 7 -41
<< metal2 >>
rect 2 -41 5 90
rect 35 46 46 49
rect 33 22 38 25
rect 35 -17 38 22
rect 35 -20 49 -17
<< m123contact >>
rect -8 -12 -3 -7
rect 72 -10 77 -5
<< metal3 >>
rect -3 -10 72 -7
use nand  nand_0
timestamp 1618580231
transform 1 0 77 0 1 3
box 0 -35 34 27
use inv  inv_0
timestamp 1618579805
transform 1 0 43 0 1 -3
box 0 -15 24 33
use nor  nor_1
timestamp 1618580541
transform 1 0 -2 0 -1 -5
box 0 -30 34 39
use nor  nor_0
timestamp 1618580541
transform 1 0 -2 0 1 54
box 0 -30 34 39
<< labels >>
rlabel metal1 -9 49 -9 52 3 p0
<< end >>
